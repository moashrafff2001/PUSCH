module Twiddle2048 #(
    parameter   TW_FF = 0   //  Use Output Register
)(
    input           clk,  //  Master Clock
    input   [11:0]   addr,   //  Twiddle Factor Number
    output  [25:0]  tw_re,  //  Twiddle Factor (Real)
    output  [25:0]  tw_im   //  Twiddle Factor (Imag)
);

wire[25:0]  wn_re[0:2047];   //  Twiddle Table (Real)
wire[25:0]  wn_im[0:2047];   //  Twiddle Table (Imag)
wire[25:0]  mx_re;          //  Multiplexer output (Real)
wire[25:0]  mx_im;          //  Multiplexer output (Imag)
reg [25:0]  ff_re;          //  Register output (Real)
reg [25:0]  ff_im;          //  Register output (Imag)

assign  mx_re = wn_re[addr];
assign  mx_im = wn_im[addr];

always @(posedge clk) begin
    ff_re <= mx_re;
    ff_im <= mx_im;
end

assign  tw_re = TW_FF ? ff_re : mx_re;
assign  tw_im = TW_FF ? ff_im : mx_im;
assign wn_re[0] = 26'b00000000000000010000000000; assign wn_im[0] = 26'b00000000000000000000000000; 
assign wn_re[1] = 26'b00000000000000001111111111; assign wn_im[1] = 26'b11111111111111111111111100; 
assign wn_re[2] = 26'b00000000000000001111111111; assign wn_im[2] = 26'b11111111111111111111111001; 
assign wn_re[3] = 26'b00000000000000001111111111; assign wn_im[3] = 26'b11111111111111111111110110; 
assign wn_re[4] = 26'b00000000000000001111111111; assign wn_im[4] = 26'b11111111111111111111110011; 
assign wn_re[5] = 26'b00000000000000001111111111; assign wn_im[5] = 26'b11111111111111111111110000; 
assign wn_re[6] = 26'b00000000000000001111111111; assign wn_im[6] = 26'b11111111111111111111101101; 
assign wn_re[7] = 26'b00000000000000001111111111; assign wn_im[7] = 26'b11111111111111111111101010; 
assign wn_re[8] = 26'b00000000000000001111111111; assign wn_im[8] = 26'b11111111111111111111100110; 
assign wn_re[9] = 26'b00000000000000001111111111; assign wn_im[9] = 26'b11111111111111111111100011; 
assign wn_re[10] = 26'b00000000000000001111111111; assign wn_im[10] = 26'b11111111111111111111100000; 
assign wn_re[11] = 26'b00000000000000001111111111; assign wn_im[11] = 26'b11111111111111111111011101; 
assign wn_re[12] = 26'b00000000000000001111111111; assign wn_im[12] = 26'b11111111111111111111011010; 
assign wn_re[13] = 26'b00000000000000001111111111; assign wn_im[13] = 26'b11111111111111111111010111; 
assign wn_re[14] = 26'b00000000000000001111111111; assign wn_im[14] = 26'b11111111111111111111010100; 
assign wn_re[15] = 26'b00000000000000001111111110; assign wn_im[15] = 26'b11111111111111111111010000; 
assign wn_re[16] = 26'b00000000000000001111111110; assign wn_im[16] = 26'b11111111111111111111001101; 
assign wn_re[17] = 26'b00000000000000001111111110; assign wn_im[17] = 26'b11111111111111111111001010; 
assign wn_re[18] = 26'b00000000000000001111111110; assign wn_im[18] = 26'b11111111111111111111000111; 
assign wn_re[19] = 26'b00000000000000001111111110; assign wn_im[19] = 26'b11111111111111111111000100; 
assign wn_re[20] = 26'b00000000000000001111111110; assign wn_im[20] = 26'b11111111111111111111000001; 
assign wn_re[21] = 26'b00000000000000001111111101; assign wn_im[21] = 26'b11111111111111111110111110; 
assign wn_re[22] = 26'b00000000000000001111111101; assign wn_im[22] = 26'b11111111111111111110111010; 
assign wn_re[23] = 26'b00000000000000001111111101; assign wn_im[23] = 26'b11111111111111111110110111; 
assign wn_re[24] = 26'b00000000000000001111111101; assign wn_im[24] = 26'b11111111111111111110110100; 
assign wn_re[25] = 26'b00000000000000001111111100; assign wn_im[25] = 26'b11111111111111111110110001; 
assign wn_re[26] = 26'b00000000000000001111111100; assign wn_im[26] = 26'b11111111111111111110101110; 
assign wn_re[27] = 26'b00000000000000001111111100; assign wn_im[27] = 26'b11111111111111111110101011; 
assign wn_re[28] = 26'b00000000000000001111111100; assign wn_im[28] = 26'b11111111111111111110101000; 
assign wn_re[29] = 26'b00000000000000001111111011; assign wn_im[29] = 26'b11111111111111111110100101; 
assign wn_re[30] = 26'b00000000000000001111111011; assign wn_im[30] = 26'b11111111111111111110100001; 
assign wn_re[31] = 26'b00000000000000001111111011; assign wn_im[31] = 26'b11111111111111111110011110; 
assign wn_re[32] = 26'b00000000000000001111111011; assign wn_im[32] = 26'b11111111111111111110011011; 
assign wn_re[33] = 26'b00000000000000001111111010; assign wn_im[33] = 26'b11111111111111111110011000; 
assign wn_re[34] = 26'b00000000000000001111111010; assign wn_im[34] = 26'b11111111111111111110010101; 
assign wn_re[35] = 26'b00000000000000001111111010; assign wn_im[35] = 26'b11111111111111111110010010; 
assign wn_re[36] = 26'b00000000000000001111111001; assign wn_im[36] = 26'b11111111111111111110001111; 
assign wn_re[37] = 26'b00000000000000001111111001; assign wn_im[37] = 26'b11111111111111111110001100; 
assign wn_re[38] = 26'b00000000000000001111111001; assign wn_im[38] = 26'b11111111111111111110001000; 
assign wn_re[39] = 26'b00000000000000001111111000; assign wn_im[39] = 26'b11111111111111111110000101; 
assign wn_re[40] = 26'b00000000000000001111111000; assign wn_im[40] = 26'b11111111111111111110000010; 
assign wn_re[41] = 26'b00000000000000001111110111; assign wn_im[41] = 26'b11111111111111111101111111; 
assign wn_re[42] = 26'b00000000000000001111110111; assign wn_im[42] = 26'b11111111111111111101111100; 
assign wn_re[43] = 26'b00000000000000001111110111; assign wn_im[43] = 26'b11111111111111111101111001; 
assign wn_re[44] = 26'b00000000000000001111110110; assign wn_im[44] = 26'b11111111111111111101110110; 
assign wn_re[45] = 26'b00000000000000001111110110; assign wn_im[45] = 26'b11111111111111111101110011; 
assign wn_re[46] = 26'b00000000000000001111110101; assign wn_im[46] = 26'b11111111111111111101101111; 
assign wn_re[47] = 26'b00000000000000001111110101; assign wn_im[47] = 26'b11111111111111111101101100; 
assign wn_re[48] = 26'b00000000000000001111110100; assign wn_im[48] = 26'b11111111111111111101101001; 
assign wn_re[49] = 26'b00000000000000001111110100; assign wn_im[49] = 26'b11111111111111111101100110; 
assign wn_re[50] = 26'b00000000000000001111110011; assign wn_im[50] = 26'b11111111111111111101100011; 
assign wn_re[51] = 26'b00000000000000001111110011; assign wn_im[51] = 26'b11111111111111111101100000; 
assign wn_re[52] = 26'b00000000000000001111110010; assign wn_im[52] = 26'b11111111111111111101011101; 
assign wn_re[53] = 26'b00000000000000001111110010; assign wn_im[53] = 26'b11111111111111111101011010; 
assign wn_re[54] = 26'b00000000000000001111110001; assign wn_im[54] = 26'b11111111111111111101010111; 
assign wn_re[55] = 26'b00000000000000001111110001; assign wn_im[55] = 26'b11111111111111111101010100; 
assign wn_re[56] = 26'b00000000000000001111110000; assign wn_im[56] = 26'b11111111111111111101010000; 
assign wn_re[57] = 26'b00000000000000001111110000; assign wn_im[57] = 26'b11111111111111111101001101; 
assign wn_re[58] = 26'b00000000000000001111101111; assign wn_im[58] = 26'b11111111111111111101001010; 
assign wn_re[59] = 26'b00000000000000001111101111; assign wn_im[59] = 26'b11111111111111111101000111; 
assign wn_re[60] = 26'b00000000000000001111101110; assign wn_im[60] = 26'b11111111111111111101000100; 
assign wn_re[61] = 26'b00000000000000001111101110; assign wn_im[61] = 26'b11111111111111111101000001; 
assign wn_re[62] = 26'b00000000000000001111101101; assign wn_im[62] = 26'b11111111111111111100111110; 
assign wn_re[63] = 26'b00000000000000001111101100; assign wn_im[63] = 26'b11111111111111111100111011; 
assign wn_re[64] = 26'b00000000000000001111101100; assign wn_im[64] = 26'b11111111111111111100111000; 
assign wn_re[65] = 26'b00000000000000001111101011; assign wn_im[65] = 26'b11111111111111111100110101; 
assign wn_re[66] = 26'b00000000000000001111101011; assign wn_im[66] = 26'b11111111111111111100110010; 
assign wn_re[67] = 26'b00000000000000001111101010; assign wn_im[67] = 26'b11111111111111111100101110; 
assign wn_re[68] = 26'b00000000000000001111101001; assign wn_im[68] = 26'b11111111111111111100101011; 
assign wn_re[69] = 26'b00000000000000001111101001; assign wn_im[69] = 26'b11111111111111111100101000; 
assign wn_re[70] = 26'b00000000000000001111101000; assign wn_im[70] = 26'b11111111111111111100100101; 
assign wn_re[71] = 26'b00000000000000001111100111; assign wn_im[71] = 26'b11111111111111111100100010; 
assign wn_re[72] = 26'b00000000000000001111100111; assign wn_im[72] = 26'b11111111111111111100011111; 
assign wn_re[73] = 26'b00000000000000001111100110; assign wn_im[73] = 26'b11111111111111111100011100; 
assign wn_re[74] = 26'b00000000000000001111100101; assign wn_im[74] = 26'b11111111111111111100011001; 
assign wn_re[75] = 26'b00000000000000001111100101; assign wn_im[75] = 26'b11111111111111111100010110; 
assign wn_re[76] = 26'b00000000000000001111100100; assign wn_im[76] = 26'b11111111111111111100010011; 
assign wn_re[77] = 26'b00000000000000001111100011; assign wn_im[77] = 26'b11111111111111111100010000; 
assign wn_re[78] = 26'b00000000000000001111100010; assign wn_im[78] = 26'b11111111111111111100001101; 
assign wn_re[79] = 26'b00000000000000001111100010; assign wn_im[79] = 26'b11111111111111111100001010; 
assign wn_re[80] = 26'b00000000000000001111100001; assign wn_im[80] = 26'b11111111111111111100000111; 
assign wn_re[81] = 26'b00000000000000001111100000; assign wn_im[81] = 26'b11111111111111111100000100; 
assign wn_re[82] = 26'b00000000000000001111011111; assign wn_im[82] = 26'b11111111111111111100000001; 
assign wn_re[83] = 26'b00000000000000001111011110; assign wn_im[83] = 26'b11111111111111111011111110; 
assign wn_re[84] = 26'b00000000000000001111011110; assign wn_im[84] = 26'b11111111111111111011111011; 
assign wn_re[85] = 26'b00000000000000001111011101; assign wn_im[85] = 26'b11111111111111111011110111; 
assign wn_re[86] = 26'b00000000000000001111011100; assign wn_im[86] = 26'b11111111111111111011110100; 
assign wn_re[87] = 26'b00000000000000001111011011; assign wn_im[87] = 26'b11111111111111111011110001; 
assign wn_re[88] = 26'b00000000000000001111011010; assign wn_im[88] = 26'b11111111111111111011101110; 
assign wn_re[89] = 26'b00000000000000001111011010; assign wn_im[89] = 26'b11111111111111111011101011; 
assign wn_re[90] = 26'b00000000000000001111011001; assign wn_im[90] = 26'b11111111111111111011101000; 
assign wn_re[91] = 26'b00000000000000001111011000; assign wn_im[91] = 26'b11111111111111111011100101; 
assign wn_re[92] = 26'b00000000000000001111010111; assign wn_im[92] = 26'b11111111111111111011100010; 
assign wn_re[93] = 26'b00000000000000001111010110; assign wn_im[93] = 26'b11111111111111111011011111; 
assign wn_re[94] = 26'b00000000000000001111010101; assign wn_im[94] = 26'b11111111111111111011011100; 
assign wn_re[95] = 26'b00000000000000001111010100; assign wn_im[95] = 26'b11111111111111111011011001; 
assign wn_re[96] = 26'b00000000000000001111010011; assign wn_im[96] = 26'b11111111111111111011010110; 
assign wn_re[97] = 26'b00000000000000001111010010; assign wn_im[97] = 26'b11111111111111111011010011; 
assign wn_re[98] = 26'b00000000000000001111010010; assign wn_im[98] = 26'b11111111111111111011010000; 
assign wn_re[99] = 26'b00000000000000001111010001; assign wn_im[99] = 26'b11111111111111111011001101; 
assign wn_re[100] = 26'b00000000000000001111010000; assign wn_im[100] = 26'b11111111111111111011001010; 
assign wn_re[101] = 26'b00000000000000001111001111; assign wn_im[101] = 26'b11111111111111111011000111; 
assign wn_re[102] = 26'b00000000000000001111001110; assign wn_im[102] = 26'b11111111111111111011000100; 
assign wn_re[103] = 26'b00000000000000001111001101; assign wn_im[103] = 26'b11111111111111111011000001; 
assign wn_re[104] = 26'b00000000000000001111001100; assign wn_im[104] = 26'b11111111111111111010111110; 
assign wn_re[105] = 26'b00000000000000001111001011; assign wn_im[105] = 26'b11111111111111111010111011; 
assign wn_re[106] = 26'b00000000000000001111001010; assign wn_im[106] = 26'b11111111111111111010111000; 
assign wn_re[107] = 26'b00000000000000001111001001; assign wn_im[107] = 26'b11111111111111111010110101; 
assign wn_re[108] = 26'b00000000000000001111001000; assign wn_im[108] = 26'b11111111111111111010110010; 
assign wn_re[109] = 26'b00000000000000001111000111; assign wn_im[109] = 26'b11111111111111111010101111; 
assign wn_re[110] = 26'b00000000000000001111000110; assign wn_im[110] = 26'b11111111111111111010101100; 
assign wn_re[111] = 26'b00000000000000001111000101; assign wn_im[111] = 26'b11111111111111111010101001; 
assign wn_re[112] = 26'b00000000000000001111000100; assign wn_im[112] = 26'b11111111111111111010100111; 
assign wn_re[113] = 26'b00000000000000001111000011; assign wn_im[113] = 26'b11111111111111111010100100; 
assign wn_re[114] = 26'b00000000000000001111000010; assign wn_im[114] = 26'b11111111111111111010100001; 
assign wn_re[115] = 26'b00000000000000001111000000; assign wn_im[115] = 26'b11111111111111111010011110; 
assign wn_re[116] = 26'b00000000000000001110111111; assign wn_im[116] = 26'b11111111111111111010011011; 
assign wn_re[117] = 26'b00000000000000001110111110; assign wn_im[117] = 26'b11111111111111111010011000; 
assign wn_re[118] = 26'b00000000000000001110111101; assign wn_im[118] = 26'b11111111111111111010010101; 
assign wn_re[119] = 26'b00000000000000001110111100; assign wn_im[119] = 26'b11111111111111111010010010; 
assign wn_re[120] = 26'b00000000000000001110111011; assign wn_im[120] = 26'b11111111111111111010001111; 
assign wn_re[121] = 26'b00000000000000001110111010; assign wn_im[121] = 26'b11111111111111111010001100; 
assign wn_re[122] = 26'b00000000000000001110111001; assign wn_im[122] = 26'b11111111111111111010001001; 
assign wn_re[123] = 26'b00000000000000001110110111; assign wn_im[123] = 26'b11111111111111111010000110; 
assign wn_re[124] = 26'b00000000000000001110110110; assign wn_im[124] = 26'b11111111111111111010000011; 
assign wn_re[125] = 26'b00000000000000001110110101; assign wn_im[125] = 26'b11111111111111111010000000; 
assign wn_re[126] = 26'b00000000000000001110110100; assign wn_im[126] = 26'b11111111111111111001111101; 
assign wn_re[127] = 26'b00000000000000001110110011; assign wn_im[127] = 26'b11111111111111111001111011; 
assign wn_re[128] = 26'b00000000000000001110110010; assign wn_im[128] = 26'b11111111111111111001111000; 
assign wn_re[129] = 26'b00000000000000001110110000; assign wn_im[129] = 26'b11111111111111111001110101; 
assign wn_re[130] = 26'b00000000000000001110101111; assign wn_im[130] = 26'b11111111111111111001110010; 
assign wn_re[131] = 26'b00000000000000001110101110; assign wn_im[131] = 26'b11111111111111111001101111; 
assign wn_re[132] = 26'b00000000000000001110101101; assign wn_im[132] = 26'b11111111111111111001101100; 
assign wn_re[133] = 26'b00000000000000001110101011; assign wn_im[133] = 26'b11111111111111111001101001; 
assign wn_re[134] = 26'b00000000000000001110101010; assign wn_im[134] = 26'b11111111111111111001100110; 
assign wn_re[135] = 26'b00000000000000001110101001; assign wn_im[135] = 26'b11111111111111111001100011; 
assign wn_re[136] = 26'b00000000000000001110101000; assign wn_im[136] = 26'b11111111111111111001100001; 
assign wn_re[137] = 26'b00000000000000001110100110; assign wn_im[137] = 26'b11111111111111111001011110; 
assign wn_re[138] = 26'b00000000000000001110100101; assign wn_im[138] = 26'b11111111111111111001011011; 
assign wn_re[139] = 26'b00000000000000001110100100; assign wn_im[139] = 26'b11111111111111111001011000; 
assign wn_re[140] = 26'b00000000000000001110100010; assign wn_im[140] = 26'b11111111111111111001010101; 
assign wn_re[141] = 26'b00000000000000001110100001; assign wn_im[141] = 26'b11111111111111111001010010; 
assign wn_re[142] = 26'b00000000000000001110100000; assign wn_im[142] = 26'b11111111111111111001001111; 
assign wn_re[143] = 26'b00000000000000001110011111; assign wn_im[143] = 26'b11111111111111111001001101; 
assign wn_re[144] = 26'b00000000000000001110011101; assign wn_im[144] = 26'b11111111111111111001001010; 
assign wn_re[145] = 26'b00000000000000001110011100; assign wn_im[145] = 26'b11111111111111111001000111; 
assign wn_re[146] = 26'b00000000000000001110011010; assign wn_im[146] = 26'b11111111111111111001000100; 
assign wn_re[147] = 26'b00000000000000001110011001; assign wn_im[147] = 26'b11111111111111111001000001; 
assign wn_re[148] = 26'b00000000000000001110011000; assign wn_im[148] = 26'b11111111111111111000111110; 
assign wn_re[149] = 26'b00000000000000001110010110; assign wn_im[149] = 26'b11111111111111111000111100; 
assign wn_re[150] = 26'b00000000000000001110010101; assign wn_im[150] = 26'b11111111111111111000111001; 
assign wn_re[151] = 26'b00000000000000001110010100; assign wn_im[151] = 26'b11111111111111111000110110; 
assign wn_re[152] = 26'b00000000000000001110010010; assign wn_im[152] = 26'b11111111111111111000110011; 
assign wn_re[153] = 26'b00000000000000001110010001; assign wn_im[153] = 26'b11111111111111111000110000; 
assign wn_re[154] = 26'b00000000000000001110001111; assign wn_im[154] = 26'b11111111111111111000101101; 
assign wn_re[155] = 26'b00000000000000001110001110; assign wn_im[155] = 26'b11111111111111111000101011; 
assign wn_re[156] = 26'b00000000000000001110001100; assign wn_im[156] = 26'b11111111111111111000101000; 
assign wn_re[157] = 26'b00000000000000001110001011; assign wn_im[157] = 26'b11111111111111111000100101; 
assign wn_re[158] = 26'b00000000000000001110001010; assign wn_im[158] = 26'b11111111111111111000100010; 
assign wn_re[159] = 26'b00000000000000001110001000; assign wn_im[159] = 26'b11111111111111111000100000; 
assign wn_re[160] = 26'b00000000000000001110000111; assign wn_im[160] = 26'b11111111111111111000011101; 
assign wn_re[161] = 26'b00000000000000001110000101; assign wn_im[161] = 26'b11111111111111111000011010; 
assign wn_re[162] = 26'b00000000000000001110000100; assign wn_im[162] = 26'b11111111111111111000010111; 
assign wn_re[163] = 26'b00000000000000001110000010; assign wn_im[163] = 26'b11111111111111111000010100; 
assign wn_re[164] = 26'b00000000000000001110000001; assign wn_im[164] = 26'b11111111111111111000010010; 
assign wn_re[165] = 26'b00000000000000001101111111; assign wn_im[165] = 26'b11111111111111111000001111; 
assign wn_re[166] = 26'b00000000000000001101111110; assign wn_im[166] = 26'b11111111111111111000001100; 
assign wn_re[167] = 26'b00000000000000001101111100; assign wn_im[167] = 26'b11111111111111111000001010; 
assign wn_re[168] = 26'b00000000000000001101111010; assign wn_im[168] = 26'b11111111111111111000000111; 
assign wn_re[169] = 26'b00000000000000001101111001; assign wn_im[169] = 26'b11111111111111111000000100; 
assign wn_re[170] = 26'b00000000000000001101110111; assign wn_im[170] = 26'b11111111111111111000000001; 
assign wn_re[171] = 26'b00000000000000001101110110; assign wn_im[171] = 26'b11111111111111110111111111; 
assign wn_re[172] = 26'b00000000000000001101110100; assign wn_im[172] = 26'b11111111111111110111111100; 
assign wn_re[173] = 26'b00000000000000001101110011; assign wn_im[173] = 26'b11111111111111110111111001; 
assign wn_re[174] = 26'b00000000000000001101110001; assign wn_im[174] = 26'b11111111111111110111110110; 
assign wn_re[175] = 26'b00000000000000001101101111; assign wn_im[175] = 26'b11111111111111110111110100; 
assign wn_re[176] = 26'b00000000000000001101101110; assign wn_im[176] = 26'b11111111111111110111110001; 
assign wn_re[177] = 26'b00000000000000001101101100; assign wn_im[177] = 26'b11111111111111110111101110; 
assign wn_re[178] = 26'b00000000000000001101101011; assign wn_im[178] = 26'b11111111111111110111101100; 
assign wn_re[179] = 26'b00000000000000001101101001; assign wn_im[179] = 26'b11111111111111110111101001; 
assign wn_re[180] = 26'b00000000000000001101100111; assign wn_im[180] = 26'b11111111111111110111100110; 
assign wn_re[181] = 26'b00000000000000001101100110; assign wn_im[181] = 26'b11111111111111110111100100; 
assign wn_re[182] = 26'b00000000000000001101100100; assign wn_im[182] = 26'b11111111111111110111100001; 
assign wn_re[183] = 26'b00000000000000001101100010; assign wn_im[183] = 26'b11111111111111110111011110; 
assign wn_re[184] = 26'b00000000000000001101100001; assign wn_im[184] = 26'b11111111111111110111011100; 
assign wn_re[185] = 26'b00000000000000001101011111; assign wn_im[185] = 26'b11111111111111110111011001; 
assign wn_re[186] = 26'b00000000000000001101011101; assign wn_im[186] = 26'b11111111111111110111010110; 
assign wn_re[187] = 26'b00000000000000001101011100; assign wn_im[187] = 26'b11111111111111110111010100; 
assign wn_re[188] = 26'b00000000000000001101011010; assign wn_im[188] = 26'b11111111111111110111010001; 
assign wn_re[189] = 26'b00000000000000001101011000; assign wn_im[189] = 26'b11111111111111110111001110; 
assign wn_re[190] = 26'b00000000000000001101010110; assign wn_im[190] = 26'b11111111111111110111001100; 
assign wn_re[191] = 26'b00000000000000001101010101; assign wn_im[191] = 26'b11111111111111110111001001; 
assign wn_re[192] = 26'b00000000000000001101010011; assign wn_im[192] = 26'b11111111111111110111000111; 
assign wn_re[193] = 26'b00000000000000001101010001; assign wn_im[193] = 26'b11111111111111110111000100; 
assign wn_re[194] = 26'b00000000000000001101001111; assign wn_im[194] = 26'b11111111111111110111000001; 
assign wn_re[195] = 26'b00000000000000001101001110; assign wn_im[195] = 26'b11111111111111110110111111; 
assign wn_re[196] = 26'b00000000000000001101001100; assign wn_im[196] = 26'b11111111111111110110111100; 
assign wn_re[197] = 26'b00000000000000001101001010; assign wn_im[197] = 26'b11111111111111110110111010; 
assign wn_re[198] = 26'b00000000000000001101001000; assign wn_im[198] = 26'b11111111111111110110110111; 
assign wn_re[199] = 26'b00000000000000001101000111; assign wn_im[199] = 26'b11111111111111110110110100; 
assign wn_re[200] = 26'b00000000000000001101000101; assign wn_im[200] = 26'b11111111111111110110110010; 
assign wn_re[201] = 26'b00000000000000001101000011; assign wn_im[201] = 26'b11111111111111110110101111; 
assign wn_re[202] = 26'b00000000000000001101000001; assign wn_im[202] = 26'b11111111111111110110101101; 
assign wn_re[203] = 26'b00000000000000001100111111; assign wn_im[203] = 26'b11111111111111110110101010; 
assign wn_re[204] = 26'b00000000000000001100111101; assign wn_im[204] = 26'b11111111111111110110101000; 
assign wn_re[205] = 26'b00000000000000001100111100; assign wn_im[205] = 26'b11111111111111110110100101; 
assign wn_re[206] = 26'b00000000000000001100111010; assign wn_im[206] = 26'b11111111111111110110100011; 
assign wn_re[207] = 26'b00000000000000001100111000; assign wn_im[207] = 26'b11111111111111110110100000; 
assign wn_re[208] = 26'b00000000000000001100110110; assign wn_im[208] = 26'b11111111111111110110011110; 
assign wn_re[209] = 26'b00000000000000001100110100; assign wn_im[209] = 26'b11111111111111110110011011; 
assign wn_re[210] = 26'b00000000000000001100110010; assign wn_im[210] = 26'b11111111111111110110011000; 
assign wn_re[211] = 26'b00000000000000001100110000; assign wn_im[211] = 26'b11111111111111110110010110; 
assign wn_re[212] = 26'b00000000000000001100101110; assign wn_im[212] = 26'b11111111111111110110010011; 
assign wn_re[213] = 26'b00000000000000001100101101; assign wn_im[213] = 26'b11111111111111110110010001; 
assign wn_re[214] = 26'b00000000000000001100101011; assign wn_im[214] = 26'b11111111111111110110001110; 
assign wn_re[215] = 26'b00000000000000001100101001; assign wn_im[215] = 26'b11111111111111110110001100; 
assign wn_re[216] = 26'b00000000000000001100100111; assign wn_im[216] = 26'b11111111111111110110001010; 
assign wn_re[217] = 26'b00000000000000001100100101; assign wn_im[217] = 26'b11111111111111110110000111; 
assign wn_re[218] = 26'b00000000000000001100100011; assign wn_im[218] = 26'b11111111111111110110000101; 
assign wn_re[219] = 26'b00000000000000001100100001; assign wn_im[219] = 26'b11111111111111110110000010; 
assign wn_re[220] = 26'b00000000000000001100011111; assign wn_im[220] = 26'b11111111111111110110000000; 
assign wn_re[221] = 26'b00000000000000001100011101; assign wn_im[221] = 26'b11111111111111110101111101; 
assign wn_re[222] = 26'b00000000000000001100011011; assign wn_im[222] = 26'b11111111111111110101111011; 
assign wn_re[223] = 26'b00000000000000001100011001; assign wn_im[223] = 26'b11111111111111110101111000; 
assign wn_re[224] = 26'b00000000000000001100010111; assign wn_im[224] = 26'b11111111111111110101110110; 
assign wn_re[225] = 26'b00000000000000001100010101; assign wn_im[225] = 26'b11111111111111110101110011; 
assign wn_re[226] = 26'b00000000000000001100010011; assign wn_im[226] = 26'b11111111111111110101110001; 
assign wn_re[227] = 26'b00000000000000001100010001; assign wn_im[227] = 26'b11111111111111110101101111; 
assign wn_re[228] = 26'b00000000000000001100001111; assign wn_im[228] = 26'b11111111111111110101101100; 
assign wn_re[229] = 26'b00000000000000001100001101; assign wn_im[229] = 26'b11111111111111110101101010; 
assign wn_re[230] = 26'b00000000000000001100001011; assign wn_im[230] = 26'b11111111111111110101100111; 
assign wn_re[231] = 26'b00000000000000001100001001; assign wn_im[231] = 26'b11111111111111110101100101; 
assign wn_re[232] = 26'b00000000000000001100000111; assign wn_im[232] = 26'b11111111111111110101100011; 
assign wn_re[233] = 26'b00000000000000001100000101; assign wn_im[233] = 26'b11111111111111110101100000; 
assign wn_re[234] = 26'b00000000000000001100000011; assign wn_im[234] = 26'b11111111111111110101011110; 
assign wn_re[235] = 26'b00000000000000001100000001; assign wn_im[235] = 26'b11111111111111110101011100; 
assign wn_re[236] = 26'b00000000000000001011111111; assign wn_im[236] = 26'b11111111111111110101011001; 
assign wn_re[237] = 26'b00000000000000001011111101; assign wn_im[237] = 26'b11111111111111110101010111; 
assign wn_re[238] = 26'b00000000000000001011111010; assign wn_im[238] = 26'b11111111111111110101010100; 
assign wn_re[239] = 26'b00000000000000001011111000; assign wn_im[239] = 26'b11111111111111110101010010; 
assign wn_re[240] = 26'b00000000000000001011110110; assign wn_im[240] = 26'b11111111111111110101010000; 
assign wn_re[241] = 26'b00000000000000001011110100; assign wn_im[241] = 26'b11111111111111110101001101; 
assign wn_re[242] = 26'b00000000000000001011110010; assign wn_im[242] = 26'b11111111111111110101001011; 
assign wn_re[243] = 26'b00000000000000001011110000; assign wn_im[243] = 26'b11111111111111110101001001; 
assign wn_re[244] = 26'b00000000000000001011101110; assign wn_im[244] = 26'b11111111111111110101000111; 
assign wn_re[245] = 26'b00000000000000001011101100; assign wn_im[245] = 26'b11111111111111110101000100; 
assign wn_re[246] = 26'b00000000000000001011101001; assign wn_im[246] = 26'b11111111111111110101000010; 
assign wn_re[247] = 26'b00000000000000001011100111; assign wn_im[247] = 26'b11111111111111110101000000; 
assign wn_re[248] = 26'b00000000000000001011100101; assign wn_im[248] = 26'b11111111111111110100111101; 
assign wn_re[249] = 26'b00000000000000001011100011; assign wn_im[249] = 26'b11111111111111110100111011; 
assign wn_re[250] = 26'b00000000000000001011100001; assign wn_im[250] = 26'b11111111111111110100111001; 
assign wn_re[251] = 26'b00000000000000001011011111; assign wn_im[251] = 26'b11111111111111110100110111; 
assign wn_re[252] = 26'b00000000000000001011011100; assign wn_im[252] = 26'b11111111111111110100110100; 
assign wn_re[253] = 26'b00000000000000001011011010; assign wn_im[253] = 26'b11111111111111110100110010; 
assign wn_re[254] = 26'b00000000000000001011011000; assign wn_im[254] = 26'b11111111111111110100110000; 
assign wn_re[255] = 26'b00000000000000001011010110; assign wn_im[255] = 26'b11111111111111110100101110; 
assign wn_re[256] = 26'b00000000000000001011010100; assign wn_im[256] = 26'b11111111111111110100101011; 
assign wn_re[257] = 26'b00000000000000001011010001; assign wn_im[257] = 26'b11111111111111110100101001; 
assign wn_re[258] = 26'b00000000000000001011001111; assign wn_im[258] = 26'b11111111111111110100100111; 
assign wn_re[259] = 26'b00000000000000001011001101; assign wn_im[259] = 26'b11111111111111110100100101; 
assign wn_re[260] = 26'b00000000000000001011001011; assign wn_im[260] = 26'b11111111111111110100100011; 
assign wn_re[261] = 26'b00000000000000001011001000; assign wn_im[261] = 26'b11111111111111110100100000; 
assign wn_re[262] = 26'b00000000000000001011000110; assign wn_im[262] = 26'b11111111111111110100011110; 
assign wn_re[263] = 26'b00000000000000001011000100; assign wn_im[263] = 26'b11111111111111110100011100; 
assign wn_re[264] = 26'b00000000000000001011000010; assign wn_im[264] = 26'b11111111111111110100011010; 
assign wn_re[265] = 26'b00000000000000001010111111; assign wn_im[265] = 26'b11111111111111110100011000; 
assign wn_re[266] = 26'b00000000000000001010111101; assign wn_im[266] = 26'b11111111111111110100010110; 
assign wn_re[267] = 26'b00000000000000001010111011; assign wn_im[267] = 26'b11111111111111110100010011; 
assign wn_re[268] = 26'b00000000000000001010111000; assign wn_im[268] = 26'b11111111111111110100010001; 
assign wn_re[269] = 26'b00000000000000001010110110; assign wn_im[269] = 26'b11111111111111110100001111; 
assign wn_re[270] = 26'b00000000000000001010110100; assign wn_im[270] = 26'b11111111111111110100001101; 
assign wn_re[271] = 26'b00000000000000001010110010; assign wn_im[271] = 26'b11111111111111110100001011; 
assign wn_re[272] = 26'b00000000000000001010101111; assign wn_im[272] = 26'b11111111111111110100001001; 
assign wn_re[273] = 26'b00000000000000001010101101; assign wn_im[273] = 26'b11111111111111110100000111; 
assign wn_re[274] = 26'b00000000000000001010101011; assign wn_im[274] = 26'b11111111111111110100000101; 
assign wn_re[275] = 26'b00000000000000001010101000; assign wn_im[275] = 26'b11111111111111110100000010; 
assign wn_re[276] = 26'b00000000000000001010100110; assign wn_im[276] = 26'b11111111111111110100000000; 
assign wn_re[277] = 26'b00000000000000001010100011; assign wn_im[277] = 26'b11111111111111110011111110; 
assign wn_re[278] = 26'b00000000000000001010100001; assign wn_im[278] = 26'b11111111111111110011111100; 
assign wn_re[279] = 26'b00000000000000001010011111; assign wn_im[279] = 26'b11111111111111110011111010; 
assign wn_re[280] = 26'b00000000000000001010011100; assign wn_im[280] = 26'b11111111111111110011111000; 
assign wn_re[281] = 26'b00000000000000001010011010; assign wn_im[281] = 26'b11111111111111110011110110; 
assign wn_re[282] = 26'b00000000000000001010011000; assign wn_im[282] = 26'b11111111111111110011110100; 
assign wn_re[283] = 26'b00000000000000001010010101; assign wn_im[283] = 26'b11111111111111110011110010; 
assign wn_re[284] = 26'b00000000000000001010010011; assign wn_im[284] = 26'b11111111111111110011110000; 
assign wn_re[285] = 26'b00000000000000001010010000; assign wn_im[285] = 26'b11111111111111110011101110; 
assign wn_re[286] = 26'b00000000000000001010001110; assign wn_im[286] = 26'b11111111111111110011101100; 
assign wn_re[287] = 26'b00000000000000001010001100; assign wn_im[287] = 26'b11111111111111110011101010; 
assign wn_re[288] = 26'b00000000000000001010001001; assign wn_im[288] = 26'b11111111111111110011101000; 
assign wn_re[289] = 26'b00000000000000001010000111; assign wn_im[289] = 26'b11111111111111110011100110; 
assign wn_re[290] = 26'b00000000000000001010000100; assign wn_im[290] = 26'b11111111111111110011100100; 
assign wn_re[291] = 26'b00000000000000001010000010; assign wn_im[291] = 26'b11111111111111110011100010; 
assign wn_re[292] = 26'b00000000000000001001111111; assign wn_im[292] = 26'b11111111111111110011100000; 
assign wn_re[293] = 26'b00000000000000001001111101; assign wn_im[293] = 26'b11111111111111110011011110; 
assign wn_re[294] = 26'b00000000000000001001111010; assign wn_im[294] = 26'b11111111111111110011011100; 
assign wn_re[295] = 26'b00000000000000001001111000; assign wn_im[295] = 26'b11111111111111110011011010; 
assign wn_re[296] = 26'b00000000000000001001110101; assign wn_im[296] = 26'b11111111111111110011011000; 
assign wn_re[297] = 26'b00000000000000001001110011; assign wn_im[297] = 26'b11111111111111110011010110; 
assign wn_re[298] = 26'b00000000000000001001110001; assign wn_im[298] = 26'b11111111111111110011010100; 
assign wn_re[299] = 26'b00000000000000001001101110; assign wn_im[299] = 26'b11111111111111110011010010; 
assign wn_re[300] = 26'b00000000000000001001101100; assign wn_im[300] = 26'b11111111111111110011010001; 
assign wn_re[301] = 26'b00000000000000001001101001; assign wn_im[301] = 26'b11111111111111110011001111; 
assign wn_re[302] = 26'b00000000000000001001100111; assign wn_im[302] = 26'b11111111111111110011001101; 
assign wn_re[303] = 26'b00000000000000001001100100; assign wn_im[303] = 26'b11111111111111110011001011; 
assign wn_re[304] = 26'b00000000000000001001100001; assign wn_im[304] = 26'b11111111111111110011001001; 
assign wn_re[305] = 26'b00000000000000001001011111; assign wn_im[305] = 26'b11111111111111110011000111; 
assign wn_re[306] = 26'b00000000000000001001011100; assign wn_im[306] = 26'b11111111111111110011000101; 
assign wn_re[307] = 26'b00000000000000001001011010; assign wn_im[307] = 26'b11111111111111110011000011; 
assign wn_re[308] = 26'b00000000000000001001010111; assign wn_im[308] = 26'b11111111111111110011000010; 
assign wn_re[309] = 26'b00000000000000001001010101; assign wn_im[309] = 26'b11111111111111110011000000; 
assign wn_re[310] = 26'b00000000000000001001010010; assign wn_im[310] = 26'b11111111111111110010111110; 
assign wn_re[311] = 26'b00000000000000001001010000; assign wn_im[311] = 26'b11111111111111110010111100; 
assign wn_re[312] = 26'b00000000000000001001001101; assign wn_im[312] = 26'b11111111111111110010111010; 
assign wn_re[313] = 26'b00000000000000001001001011; assign wn_im[313] = 26'b11111111111111110010111000; 
assign wn_re[314] = 26'b00000000000000001001001000; assign wn_im[314] = 26'b11111111111111110010110111; 
assign wn_re[315] = 26'b00000000000000001001000101; assign wn_im[315] = 26'b11111111111111110010110101; 
assign wn_re[316] = 26'b00000000000000001001000011; assign wn_im[316] = 26'b11111111111111110010110011; 
assign wn_re[317] = 26'b00000000000000001001000000; assign wn_im[317] = 26'b11111111111111110010110001; 
assign wn_re[318] = 26'b00000000000000001000111110; assign wn_im[318] = 26'b11111111111111110010110000; 
assign wn_re[319] = 26'b00000000000000001000111011; assign wn_im[319] = 26'b11111111111111110010101110; 
assign wn_re[320] = 26'b00000000000000001000111000; assign wn_im[320] = 26'b11111111111111110010101100; 
assign wn_re[321] = 26'b00000000000000001000110110; assign wn_im[321] = 26'b11111111111111110010101010; 
assign wn_re[322] = 26'b00000000000000001000110011; assign wn_im[322] = 26'b11111111111111110010101001; 
assign wn_re[323] = 26'b00000000000000001000110001; assign wn_im[323] = 26'b11111111111111110010100111; 
assign wn_re[324] = 26'b00000000000000001000101110; assign wn_im[324] = 26'b11111111111111110010100101; 
assign wn_re[325] = 26'b00000000000000001000101011; assign wn_im[325] = 26'b11111111111111110010100011; 
assign wn_re[326] = 26'b00000000000000001000101001; assign wn_im[326] = 26'b11111111111111110010100010; 
assign wn_re[327] = 26'b00000000000000001000100110; assign wn_im[327] = 26'b11111111111111110010100000; 
assign wn_re[328] = 26'b00000000000000001000100011; assign wn_im[328] = 26'b11111111111111110010011110; 
assign wn_re[329] = 26'b00000000000000001000100001; assign wn_im[329] = 26'b11111111111111110010011101; 
assign wn_re[330] = 26'b00000000000000001000011110; assign wn_im[330] = 26'b11111111111111110010011011; 
assign wn_re[331] = 26'b00000000000000001000011011; assign wn_im[331] = 26'b11111111111111110010011001; 
assign wn_re[332] = 26'b00000000000000001000011001; assign wn_im[332] = 26'b11111111111111110010011000; 
assign wn_re[333] = 26'b00000000000000001000010110; assign wn_im[333] = 26'b11111111111111110010010110; 
assign wn_re[334] = 26'b00000000000000001000010011; assign wn_im[334] = 26'b11111111111111110010010100; 
assign wn_re[335] = 26'b00000000000000001000010001; assign wn_im[335] = 26'b11111111111111110010010011; 
assign wn_re[336] = 26'b00000000000000001000001110; assign wn_im[336] = 26'b11111111111111110010010001; 
assign wn_re[337] = 26'b00000000000000001000001011; assign wn_im[337] = 26'b11111111111111110010010000; 
assign wn_re[338] = 26'b00000000000000001000001001; assign wn_im[338] = 26'b11111111111111110010001110; 
assign wn_re[339] = 26'b00000000000000001000000110; assign wn_im[339] = 26'b11111111111111110010001100; 
assign wn_re[340] = 26'b00000000000000001000000011; assign wn_im[340] = 26'b11111111111111110010001011; 
assign wn_re[341] = 26'b00000000000000001000000000; assign wn_im[341] = 26'b11111111111111110010001001; 
assign wn_re[342] = 26'b00000000000000000111111110; assign wn_im[342] = 26'b11111111111111110010001000; 
assign wn_re[343] = 26'b00000000000000000111111011; assign wn_im[343] = 26'b11111111111111110010000110; 
assign wn_re[344] = 26'b00000000000000000111111000; assign wn_im[344] = 26'b11111111111111110010000101; 
assign wn_re[345] = 26'b00000000000000000111110101; assign wn_im[345] = 26'b11111111111111110010000011; 
assign wn_re[346] = 26'b00000000000000000111110011; assign wn_im[346] = 26'b11111111111111110010000001; 
assign wn_re[347] = 26'b00000000000000000111110000; assign wn_im[347] = 26'b11111111111111110010000000; 
assign wn_re[348] = 26'b00000000000000000111101101; assign wn_im[348] = 26'b11111111111111110001111110; 
assign wn_re[349] = 26'b00000000000000000111101011; assign wn_im[349] = 26'b11111111111111110001111101; 
assign wn_re[350] = 26'b00000000000000000111101000; assign wn_im[350] = 26'b11111111111111110001111011; 
assign wn_re[351] = 26'b00000000000000000111100101; assign wn_im[351] = 26'b11111111111111110001111010; 
assign wn_re[352] = 26'b00000000000000000111100010; assign wn_im[352] = 26'b11111111111111110001111000; 
assign wn_re[353] = 26'b00000000000000000111011111; assign wn_im[353] = 26'b11111111111111110001110111; 
assign wn_re[354] = 26'b00000000000000000111011101; assign wn_im[354] = 26'b11111111111111110001110101; 
assign wn_re[355] = 26'b00000000000000000111011010; assign wn_im[355] = 26'b11111111111111110001110100; 
assign wn_re[356] = 26'b00000000000000000111010111; assign wn_im[356] = 26'b11111111111111110001110011; 
assign wn_re[357] = 26'b00000000000000000111010100; assign wn_im[357] = 26'b11111111111111110001110001; 
assign wn_re[358] = 26'b00000000000000000111010010; assign wn_im[358] = 26'b11111111111111110001110000; 
assign wn_re[359] = 26'b00000000000000000111001111; assign wn_im[359] = 26'b11111111111111110001101110; 
assign wn_re[360] = 26'b00000000000000000111001100; assign wn_im[360] = 26'b11111111111111110001101101; 
assign wn_re[361] = 26'b00000000000000000111001001; assign wn_im[361] = 26'b11111111111111110001101011; 
assign wn_re[362] = 26'b00000000000000000111000110; assign wn_im[362] = 26'b11111111111111110001101010; 
assign wn_re[363] = 26'b00000000000000000111000011; assign wn_im[363] = 26'b11111111111111110001101001; 
assign wn_re[364] = 26'b00000000000000000111000001; assign wn_im[364] = 26'b11111111111111110001100111; 
assign wn_re[365] = 26'b00000000000000000110111110; assign wn_im[365] = 26'b11111111111111110001100110; 
assign wn_re[366] = 26'b00000000000000000110111011; assign wn_im[366] = 26'b11111111111111110001100101; 
assign wn_re[367] = 26'b00000000000000000110111000; assign wn_im[367] = 26'b11111111111111110001100011; 
assign wn_re[368] = 26'b00000000000000000110110101; assign wn_im[368] = 26'b11111111111111110001100010; 
assign wn_re[369] = 26'b00000000000000000110110010; assign wn_im[369] = 26'b11111111111111110001100000; 
assign wn_re[370] = 26'b00000000000000000110110000; assign wn_im[370] = 26'b11111111111111110001011111; 
assign wn_re[371] = 26'b00000000000000000110101101; assign wn_im[371] = 26'b11111111111111110001011110; 
assign wn_re[372] = 26'b00000000000000000110101010; assign wn_im[372] = 26'b11111111111111110001011101; 
assign wn_re[373] = 26'b00000000000000000110100111; assign wn_im[373] = 26'b11111111111111110001011011; 
assign wn_re[374] = 26'b00000000000000000110100100; assign wn_im[374] = 26'b11111111111111110001011010; 
assign wn_re[375] = 26'b00000000000000000110100001; assign wn_im[375] = 26'b11111111111111110001011001; 
assign wn_re[376] = 26'b00000000000000000110011110; assign wn_im[376] = 26'b11111111111111110001010111; 
assign wn_re[377] = 26'b00000000000000000110011100; assign wn_im[377] = 26'b11111111111111110001010110; 
assign wn_re[378] = 26'b00000000000000000110011001; assign wn_im[378] = 26'b11111111111111110001010101; 
assign wn_re[379] = 26'b00000000000000000110010110; assign wn_im[379] = 26'b11111111111111110001010100; 
assign wn_re[380] = 26'b00000000000000000110010011; assign wn_im[380] = 26'b11111111111111110001010010; 
assign wn_re[381] = 26'b00000000000000000110010000; assign wn_im[381] = 26'b11111111111111110001010001; 
assign wn_re[382] = 26'b00000000000000000110001101; assign wn_im[382] = 26'b11111111111111110001010000; 
assign wn_re[383] = 26'b00000000000000000110001010; assign wn_im[383] = 26'b11111111111111110001001111; 
assign wn_re[384] = 26'b00000000000000000110000111; assign wn_im[384] = 26'b11111111111111110001001101; 
assign wn_re[385] = 26'b00000000000000000110000100; assign wn_im[385] = 26'b11111111111111110001001100; 
assign wn_re[386] = 26'b00000000000000000110000010; assign wn_im[386] = 26'b11111111111111110001001011; 
assign wn_re[387] = 26'b00000000000000000101111111; assign wn_im[387] = 26'b11111111111111110001001010; 
assign wn_re[388] = 26'b00000000000000000101111100; assign wn_im[388] = 26'b11111111111111110001001001; 
assign wn_re[389] = 26'b00000000000000000101111001; assign wn_im[389] = 26'b11111111111111110001001000; 
assign wn_re[390] = 26'b00000000000000000101110110; assign wn_im[390] = 26'b11111111111111110001000110; 
assign wn_re[391] = 26'b00000000000000000101110011; assign wn_im[391] = 26'b11111111111111110001000101; 
assign wn_re[392] = 26'b00000000000000000101110000; assign wn_im[392] = 26'b11111111111111110001000100; 
assign wn_re[393] = 26'b00000000000000000101101101; assign wn_im[393] = 26'b11111111111111110001000011; 
assign wn_re[394] = 26'b00000000000000000101101010; assign wn_im[394] = 26'b11111111111111110001000010; 
assign wn_re[395] = 26'b00000000000000000101100111; assign wn_im[395] = 26'b11111111111111110001000001; 
assign wn_re[396] = 26'b00000000000000000101100100; assign wn_im[396] = 26'b11111111111111110001000000; 
assign wn_re[397] = 26'b00000000000000000101100001; assign wn_im[397] = 26'b11111111111111110000111111; 
assign wn_re[398] = 26'b00000000000000000101011110; assign wn_im[398] = 26'b11111111111111110000111101; 
assign wn_re[399] = 26'b00000000000000000101011011; assign wn_im[399] = 26'b11111111111111110000111100; 
assign wn_re[400] = 26'b00000000000000000101011000; assign wn_im[400] = 26'b11111111111111110000111011; 
assign wn_re[401] = 26'b00000000000000000101010110; assign wn_im[401] = 26'b11111111111111110000111010; 
assign wn_re[402] = 26'b00000000000000000101010011; assign wn_im[402] = 26'b11111111111111110000111001; 
assign wn_re[403] = 26'b00000000000000000101010000; assign wn_im[403] = 26'b11111111111111110000111000; 
assign wn_re[404] = 26'b00000000000000000101001101; assign wn_im[404] = 26'b11111111111111110000110111; 
assign wn_re[405] = 26'b00000000000000000101001010; assign wn_im[405] = 26'b11111111111111110000110110; 
assign wn_re[406] = 26'b00000000000000000101000111; assign wn_im[406] = 26'b11111111111111110000110101; 
assign wn_re[407] = 26'b00000000000000000101000100; assign wn_im[407] = 26'b11111111111111110000110100; 
assign wn_re[408] = 26'b00000000000000000101000001; assign wn_im[408] = 26'b11111111111111110000110011; 
assign wn_re[409] = 26'b00000000000000000100111110; assign wn_im[409] = 26'b11111111111111110000110010; 
assign wn_re[410] = 26'b00000000000000000100111011; assign wn_im[410] = 26'b11111111111111110000110001; 
assign wn_re[411] = 26'b00000000000000000100111000; assign wn_im[411] = 26'b11111111111111110000110000; 
assign wn_re[412] = 26'b00000000000000000100110101; assign wn_im[412] = 26'b11111111111111110000101111; 
assign wn_re[413] = 26'b00000000000000000100110010; assign wn_im[413] = 26'b11111111111111110000101110; 
assign wn_re[414] = 26'b00000000000000000100101111; assign wn_im[414] = 26'b11111111111111110000101101; 
assign wn_re[415] = 26'b00000000000000000100101100; assign wn_im[415] = 26'b11111111111111110000101101; 
assign wn_re[416] = 26'b00000000000000000100101001; assign wn_im[416] = 26'b11111111111111110000101100; 
assign wn_re[417] = 26'b00000000000000000100100110; assign wn_im[417] = 26'b11111111111111110000101011; 
assign wn_re[418] = 26'b00000000000000000100100011; assign wn_im[418] = 26'b11111111111111110000101010; 
assign wn_re[419] = 26'b00000000000000000100100000; assign wn_im[419] = 26'b11111111111111110000101001; 
assign wn_re[420] = 26'b00000000000000000100011101; assign wn_im[420] = 26'b11111111111111110000101000; 
assign wn_re[421] = 26'b00000000000000000100011010; assign wn_im[421] = 26'b11111111111111110000100111; 
assign wn_re[422] = 26'b00000000000000000100010111; assign wn_im[422] = 26'b11111111111111110000100110; 
assign wn_re[423] = 26'b00000000000000000100010100; assign wn_im[423] = 26'b11111111111111110000100101; 
assign wn_re[424] = 26'b00000000000000000100010001; assign wn_im[424] = 26'b11111111111111110000100101; 
assign wn_re[425] = 26'b00000000000000000100001110; assign wn_im[425] = 26'b11111111111111110000100100; 
assign wn_re[426] = 26'b00000000000000000100001011; assign wn_im[426] = 26'b11111111111111110000100011; 
assign wn_re[427] = 26'b00000000000000000100001000; assign wn_im[427] = 26'b11111111111111110000100010; 
assign wn_re[428] = 26'b00000000000000000100000100; assign wn_im[428] = 26'b11111111111111110000100001; 
assign wn_re[429] = 26'b00000000000000000100000001; assign wn_im[429] = 26'b11111111111111110000100001; 
assign wn_re[430] = 26'b00000000000000000011111110; assign wn_im[430] = 26'b11111111111111110000100000; 
assign wn_re[431] = 26'b00000000000000000011111011; assign wn_im[431] = 26'b11111111111111110000011111; 
assign wn_re[432] = 26'b00000000000000000011111000; assign wn_im[432] = 26'b11111111111111110000011110; 
assign wn_re[433] = 26'b00000000000000000011110101; assign wn_im[433] = 26'b11111111111111110000011101; 
assign wn_re[434] = 26'b00000000000000000011110010; assign wn_im[434] = 26'b11111111111111110000011101; 
assign wn_re[435] = 26'b00000000000000000011101111; assign wn_im[435] = 26'b11111111111111110000011100; 
assign wn_re[436] = 26'b00000000000000000011101100; assign wn_im[436] = 26'b11111111111111110000011011; 
assign wn_re[437] = 26'b00000000000000000011101001; assign wn_im[437] = 26'b11111111111111110000011010; 
assign wn_re[438] = 26'b00000000000000000011100110; assign wn_im[438] = 26'b11111111111111110000011010; 
assign wn_re[439] = 26'b00000000000000000011100011; assign wn_im[439] = 26'b11111111111111110000011001; 
assign wn_re[440] = 26'b00000000000000000011100000; assign wn_im[440] = 26'b11111111111111110000011000; 
assign wn_re[441] = 26'b00000000000000000011011101; assign wn_im[441] = 26'b11111111111111110000011000; 
assign wn_re[442] = 26'b00000000000000000011011010; assign wn_im[442] = 26'b11111111111111110000010111; 
assign wn_re[443] = 26'b00000000000000000011010111; assign wn_im[443] = 26'b11111111111111110000010110; 
assign wn_re[444] = 26'b00000000000000000011010100; assign wn_im[444] = 26'b11111111111111110000010110; 
assign wn_re[445] = 26'b00000000000000000011010001; assign wn_im[445] = 26'b11111111111111110000010101; 
assign wn_re[446] = 26'b00000000000000000011001101; assign wn_im[446] = 26'b11111111111111110000010100; 
assign wn_re[447] = 26'b00000000000000000011001010; assign wn_im[447] = 26'b11111111111111110000010100; 
assign wn_re[448] = 26'b00000000000000000011000111; assign wn_im[448] = 26'b11111111111111110000010011; 
assign wn_re[449] = 26'b00000000000000000011000100; assign wn_im[449] = 26'b11111111111111110000010011; 
assign wn_re[450] = 26'b00000000000000000011000001; assign wn_im[450] = 26'b11111111111111110000010010; 
assign wn_re[451] = 26'b00000000000000000010111110; assign wn_im[451] = 26'b11111111111111110000010001; 
assign wn_re[452] = 26'b00000000000000000010111011; assign wn_im[452] = 26'b11111111111111110000010001; 
assign wn_re[453] = 26'b00000000000000000010111000; assign wn_im[453] = 26'b11111111111111110000010000; 
assign wn_re[454] = 26'b00000000000000000010110101; assign wn_im[454] = 26'b11111111111111110000010000; 
assign wn_re[455] = 26'b00000000000000000010110010; assign wn_im[455] = 26'b11111111111111110000001111; 
assign wn_re[456] = 26'b00000000000000000010101111; assign wn_im[456] = 26'b11111111111111110000001111; 
assign wn_re[457] = 26'b00000000000000000010101011; assign wn_im[457] = 26'b11111111111111110000001110; 
assign wn_re[458] = 26'b00000000000000000010101000; assign wn_im[458] = 26'b11111111111111110000001110; 
assign wn_re[459] = 26'b00000000000000000010100101; assign wn_im[459] = 26'b11111111111111110000001101; 
assign wn_re[460] = 26'b00000000000000000010100010; assign wn_im[460] = 26'b11111111111111110000001101; 
assign wn_re[461] = 26'b00000000000000000010011111; assign wn_im[461] = 26'b11111111111111110000001100; 
assign wn_re[462] = 26'b00000000000000000010011100; assign wn_im[462] = 26'b11111111111111110000001100; 
assign wn_re[463] = 26'b00000000000000000010011001; assign wn_im[463] = 26'b11111111111111110000001011; 
assign wn_re[464] = 26'b00000000000000000010010110; assign wn_im[464] = 26'b11111111111111110000001011; 
assign wn_re[465] = 26'b00000000000000000010010011; assign wn_im[465] = 26'b11111111111111110000001010; 
assign wn_re[466] = 26'b00000000000000000010010000; assign wn_im[466] = 26'b11111111111111110000001010; 
assign wn_re[467] = 26'b00000000000000000010001100; assign wn_im[467] = 26'b11111111111111110000001001; 
assign wn_re[468] = 26'b00000000000000000010001001; assign wn_im[468] = 26'b11111111111111110000001001; 
assign wn_re[469] = 26'b00000000000000000010000110; assign wn_im[469] = 26'b11111111111111110000001000; 
assign wn_re[470] = 26'b00000000000000000010000011; assign wn_im[470] = 26'b11111111111111110000001000; 
assign wn_re[471] = 26'b00000000000000000010000000; assign wn_im[471] = 26'b11111111111111110000001000; 
assign wn_re[472] = 26'b00000000000000000001111101; assign wn_im[472] = 26'b11111111111111110000000111; 
assign wn_re[473] = 26'b00000000000000000001111010; assign wn_im[473] = 26'b11111111111111110000000111; 
assign wn_re[474] = 26'b00000000000000000001110111; assign wn_im[474] = 26'b11111111111111110000000110; 
assign wn_re[475] = 26'b00000000000000000001110011; assign wn_im[475] = 26'b11111111111111110000000110; 
assign wn_re[476] = 26'b00000000000000000001110000; assign wn_im[476] = 26'b11111111111111110000000110; 
assign wn_re[477] = 26'b00000000000000000001101101; assign wn_im[477] = 26'b11111111111111110000000101; 
assign wn_re[478] = 26'b00000000000000000001101010; assign wn_im[478] = 26'b11111111111111110000000101; 
assign wn_re[479] = 26'b00000000000000000001100111; assign wn_im[479] = 26'b11111111111111110000000101; 
assign wn_re[480] = 26'b00000000000000000001100100; assign wn_im[480] = 26'b11111111111111110000000100; 
assign wn_re[481] = 26'b00000000000000000001100001; assign wn_im[481] = 26'b11111111111111110000000100; 
assign wn_re[482] = 26'b00000000000000000001011110; assign wn_im[482] = 26'b11111111111111110000000100; 
assign wn_re[483] = 26'b00000000000000000001011010; assign wn_im[483] = 26'b11111111111111110000000100; 
assign wn_re[484] = 26'b00000000000000000001010111; assign wn_im[484] = 26'b11111111111111110000000011; 
assign wn_re[485] = 26'b00000000000000000001010100; assign wn_im[485] = 26'b11111111111111110000000011; 
assign wn_re[486] = 26'b00000000000000000001010001; assign wn_im[486] = 26'b11111111111111110000000011; 
assign wn_re[487] = 26'b00000000000000000001001110; assign wn_im[487] = 26'b11111111111111110000000011; 
assign wn_re[488] = 26'b00000000000000000001001011; assign wn_im[488] = 26'b11111111111111110000000010; 
assign wn_re[489] = 26'b00000000000000000001001000; assign wn_im[489] = 26'b11111111111111110000000010; 
assign wn_re[490] = 26'b00000000000000000001000101; assign wn_im[490] = 26'b11111111111111110000000010; 
assign wn_re[491] = 26'b00000000000000000001000001; assign wn_im[491] = 26'b11111111111111110000000010; 
assign wn_re[492] = 26'b00000000000000000000111110; assign wn_im[492] = 26'b11111111111111110000000001; 
assign wn_re[493] = 26'b00000000000000000000111011; assign wn_im[493] = 26'b11111111111111110000000001; 
assign wn_re[494] = 26'b00000000000000000000111000; assign wn_im[494] = 26'b11111111111111110000000001; 
assign wn_re[495] = 26'b00000000000000000000110101; assign wn_im[495] = 26'b11111111111111110000000001; 
assign wn_re[496] = 26'b00000000000000000000110010; assign wn_im[496] = 26'b11111111111111110000000001; 
assign wn_re[497] = 26'b00000000000000000000101111; assign wn_im[497] = 26'b11111111111111110000000001; 
assign wn_re[498] = 26'b00000000000000000000101011; assign wn_im[498] = 26'b11111111111111110000000000; 
assign wn_re[499] = 26'b00000000000000000000101000; assign wn_im[499] = 26'b11111111111111110000000000; 
assign wn_re[500] = 26'b00000000000000000000100101; assign wn_im[500] = 26'b11111111111111110000000000; 
assign wn_re[501] = 26'b00000000000000000000100010; assign wn_im[501] = 26'b11111111111111110000000000; 
assign wn_re[502] = 26'b00000000000000000000011111; assign wn_im[502] = 26'b11111111111111110000000000; 
assign wn_re[503] = 26'b00000000000000000000011100; assign wn_im[503] = 26'b11111111111111110000000000; 
assign wn_re[504] = 26'b00000000000000000000011001; assign wn_im[504] = 26'b11111111111111110000000000; 
assign wn_re[505] = 26'b00000000000000000000010101; assign wn_im[505] = 26'b11111111111111110000000000; 
assign wn_re[506] = 26'b00000000000000000000010010; assign wn_im[506] = 26'b11111111111111110000000000; 
assign wn_re[507] = 26'b00000000000000000000001111; assign wn_im[507] = 26'b11111111111111110000000000; 
assign wn_re[508] = 26'b00000000000000000000001100; assign wn_im[508] = 26'b11111111111111110000000000; 
assign wn_re[509] = 26'b00000000000000000000001001; assign wn_im[509] = 26'b11111111111111110000000000; 
assign wn_re[510] = 26'b00000000000000000000000110; assign wn_im[510] = 26'b11111111111111110000000000; 
assign wn_re[511] = 26'b00000000000000000000000011; assign wn_im[511] = 26'b11111111111111110000000000; 
assign wn_re[512] = 26'b00000000000000000000000000; assign wn_im[512] = 26'b11111111111111110000000000; 
assign wn_re[513] = 26'b11111111111111111111111100; assign wn_im[513] = 26'b11111111111111110000000000; 
assign wn_re[514] = 26'b11111111111111111111111001; assign wn_im[514] = 26'b11111111111111110000000000; 
assign wn_re[515] = 26'b11111111111111111111110110; assign wn_im[515] = 26'b11111111111111110000000000; 
assign wn_re[516] = 26'b11111111111111111111110011; assign wn_im[516] = 26'b11111111111111110000000000; 
assign wn_re[517] = 26'b11111111111111111111110000; assign wn_im[517] = 26'b11111111111111110000000000; 
assign wn_re[518] = 26'b11111111111111111111101101; assign wn_im[518] = 26'b11111111111111110000000000; 
assign wn_re[519] = 26'b11111111111111111111101010; assign wn_im[519] = 26'b11111111111111110000000000; 
assign wn_re[520] = 26'b11111111111111111111100110; assign wn_im[520] = 26'b11111111111111110000000000; 
assign wn_re[521] = 26'b11111111111111111111100011; assign wn_im[521] = 26'b11111111111111110000000000; 
assign wn_re[522] = 26'b11111111111111111111100000; assign wn_im[522] = 26'b11111111111111110000000000; 
assign wn_re[523] = 26'b11111111111111111111011101; assign wn_im[523] = 26'b11111111111111110000000000; 
assign wn_re[524] = 26'b11111111111111111111011010; assign wn_im[524] = 26'b11111111111111110000000000; 
assign wn_re[525] = 26'b11111111111111111111010111; assign wn_im[525] = 26'b11111111111111110000000000; 
assign wn_re[526] = 26'b11111111111111111111010100; assign wn_im[526] = 26'b11111111111111110000000000; 
assign wn_re[527] = 26'b11111111111111111111010000; assign wn_im[527] = 26'b11111111111111110000000001; 
assign wn_re[528] = 26'b11111111111111111111001101; assign wn_im[528] = 26'b11111111111111110000000001; 
assign wn_re[529] = 26'b11111111111111111111001010; assign wn_im[529] = 26'b11111111111111110000000001; 
assign wn_re[530] = 26'b11111111111111111111000111; assign wn_im[530] = 26'b11111111111111110000000001; 
assign wn_re[531] = 26'b11111111111111111111000100; assign wn_im[531] = 26'b11111111111111110000000001; 
assign wn_re[532] = 26'b11111111111111111111000001; assign wn_im[532] = 26'b11111111111111110000000001; 
assign wn_re[533] = 26'b11111111111111111110111110; assign wn_im[533] = 26'b11111111111111110000000010; 
assign wn_re[534] = 26'b11111111111111111110111010; assign wn_im[534] = 26'b11111111111111110000000010; 
assign wn_re[535] = 26'b11111111111111111110110111; assign wn_im[535] = 26'b11111111111111110000000010; 
assign wn_re[536] = 26'b11111111111111111110110100; assign wn_im[536] = 26'b11111111111111110000000010; 
assign wn_re[537] = 26'b11111111111111111110110001; assign wn_im[537] = 26'b11111111111111110000000011; 
assign wn_re[538] = 26'b11111111111111111110101110; assign wn_im[538] = 26'b11111111111111110000000011; 
assign wn_re[539] = 26'b11111111111111111110101011; assign wn_im[539] = 26'b11111111111111110000000011; 
assign wn_re[540] = 26'b11111111111111111110101000; assign wn_im[540] = 26'b11111111111111110000000011; 
assign wn_re[541] = 26'b11111111111111111110100101; assign wn_im[541] = 26'b11111111111111110000000100; 
assign wn_re[542] = 26'b11111111111111111110100001; assign wn_im[542] = 26'b11111111111111110000000100; 
assign wn_re[543] = 26'b11111111111111111110011110; assign wn_im[543] = 26'b11111111111111110000000100; 
assign wn_re[544] = 26'b11111111111111111110011011; assign wn_im[544] = 26'b11111111111111110000000100; 
assign wn_re[545] = 26'b11111111111111111110011000; assign wn_im[545] = 26'b11111111111111110000000101; 
assign wn_re[546] = 26'b11111111111111111110010101; assign wn_im[546] = 26'b11111111111111110000000101; 
assign wn_re[547] = 26'b11111111111111111110010010; assign wn_im[547] = 26'b11111111111111110000000101; 
assign wn_re[548] = 26'b11111111111111111110001111; assign wn_im[548] = 26'b11111111111111110000000110; 
assign wn_re[549] = 26'b11111111111111111110001100; assign wn_im[549] = 26'b11111111111111110000000110; 
assign wn_re[550] = 26'b11111111111111111110001000; assign wn_im[550] = 26'b11111111111111110000000110; 
assign wn_re[551] = 26'b11111111111111111110000101; assign wn_im[551] = 26'b11111111111111110000000111; 
assign wn_re[552] = 26'b11111111111111111110000010; assign wn_im[552] = 26'b11111111111111110000000111; 
assign wn_re[553] = 26'b11111111111111111101111111; assign wn_im[553] = 26'b11111111111111110000001000; 
assign wn_re[554] = 26'b11111111111111111101111100; assign wn_im[554] = 26'b11111111111111110000001000; 
assign wn_re[555] = 26'b11111111111111111101111001; assign wn_im[555] = 26'b11111111111111110000001000; 
assign wn_re[556] = 26'b11111111111111111101110110; assign wn_im[556] = 26'b11111111111111110000001001; 
assign wn_re[557] = 26'b11111111111111111101110011; assign wn_im[557] = 26'b11111111111111110000001001; 
assign wn_re[558] = 26'b11111111111111111101101111; assign wn_im[558] = 26'b11111111111111110000001010; 
assign wn_re[559] = 26'b11111111111111111101101100; assign wn_im[559] = 26'b11111111111111110000001010; 
assign wn_re[560] = 26'b11111111111111111101101001; assign wn_im[560] = 26'b11111111111111110000001011; 
assign wn_re[561] = 26'b11111111111111111101100110; assign wn_im[561] = 26'b11111111111111110000001011; 
assign wn_re[562] = 26'b11111111111111111101100011; assign wn_im[562] = 26'b11111111111111110000001100; 
assign wn_re[563] = 26'b11111111111111111101100000; assign wn_im[563] = 26'b11111111111111110000001100; 
assign wn_re[564] = 26'b11111111111111111101011101; assign wn_im[564] = 26'b11111111111111110000001101; 
assign wn_re[565] = 26'b11111111111111111101011010; assign wn_im[565] = 26'b11111111111111110000001101; 
assign wn_re[566] = 26'b11111111111111111101010111; assign wn_im[566] = 26'b11111111111111110000001110; 
assign wn_re[567] = 26'b11111111111111111101010100; assign wn_im[567] = 26'b11111111111111110000001110; 
assign wn_re[568] = 26'b11111111111111111101010000; assign wn_im[568] = 26'b11111111111111110000001111; 
assign wn_re[569] = 26'b11111111111111111101001101; assign wn_im[569] = 26'b11111111111111110000001111; 
assign wn_re[570] = 26'b11111111111111111101001010; assign wn_im[570] = 26'b11111111111111110000010000; 
assign wn_re[571] = 26'b11111111111111111101000111; assign wn_im[571] = 26'b11111111111111110000010000; 
assign wn_re[572] = 26'b11111111111111111101000100; assign wn_im[572] = 26'b11111111111111110000010001; 
assign wn_re[573] = 26'b11111111111111111101000001; assign wn_im[573] = 26'b11111111111111110000010001; 
assign wn_re[574] = 26'b11111111111111111100111110; assign wn_im[574] = 26'b11111111111111110000010010; 
assign wn_re[575] = 26'b11111111111111111100111011; assign wn_im[575] = 26'b11111111111111110000010011; 
assign wn_re[576] = 26'b11111111111111111100111000; assign wn_im[576] = 26'b11111111111111110000010011; 
assign wn_re[577] = 26'b11111111111111111100110101; assign wn_im[577] = 26'b11111111111111110000010100; 
assign wn_re[578] = 26'b11111111111111111100110010; assign wn_im[578] = 26'b11111111111111110000010100; 
assign wn_re[579] = 26'b11111111111111111100101110; assign wn_im[579] = 26'b11111111111111110000010101; 
assign wn_re[580] = 26'b11111111111111111100101011; assign wn_im[580] = 26'b11111111111111110000010110; 
assign wn_re[581] = 26'b11111111111111111100101000; assign wn_im[581] = 26'b11111111111111110000010110; 
assign wn_re[582] = 26'b11111111111111111100100101; assign wn_im[582] = 26'b11111111111111110000010111; 
assign wn_re[583] = 26'b11111111111111111100100010; assign wn_im[583] = 26'b11111111111111110000011000; 
assign wn_re[584] = 26'b11111111111111111100011111; assign wn_im[584] = 26'b11111111111111110000011000; 
assign wn_re[585] = 26'b11111111111111111100011100; assign wn_im[585] = 26'b11111111111111110000011001; 
assign wn_re[586] = 26'b11111111111111111100011001; assign wn_im[586] = 26'b11111111111111110000011010; 
assign wn_re[587] = 26'b11111111111111111100010110; assign wn_im[587] = 26'b11111111111111110000011010; 
assign wn_re[588] = 26'b11111111111111111100010011; assign wn_im[588] = 26'b11111111111111110000011011; 
assign wn_re[589] = 26'b11111111111111111100010000; assign wn_im[589] = 26'b11111111111111110000011100; 
assign wn_re[590] = 26'b11111111111111111100001101; assign wn_im[590] = 26'b11111111111111110000011101; 
assign wn_re[591] = 26'b11111111111111111100001010; assign wn_im[591] = 26'b11111111111111110000011101; 
assign wn_re[592] = 26'b11111111111111111100000111; assign wn_im[592] = 26'b11111111111111110000011110; 
assign wn_re[593] = 26'b11111111111111111100000100; assign wn_im[593] = 26'b11111111111111110000011111; 
assign wn_re[594] = 26'b11111111111111111100000001; assign wn_im[594] = 26'b11111111111111110000100000; 
assign wn_re[595] = 26'b11111111111111111011111110; assign wn_im[595] = 26'b11111111111111110000100001; 
assign wn_re[596] = 26'b11111111111111111011111011; assign wn_im[596] = 26'b11111111111111110000100001; 
assign wn_re[597] = 26'b11111111111111111011110111; assign wn_im[597] = 26'b11111111111111110000100010; 
assign wn_re[598] = 26'b11111111111111111011110100; assign wn_im[598] = 26'b11111111111111110000100011; 
assign wn_re[599] = 26'b11111111111111111011110001; assign wn_im[599] = 26'b11111111111111110000100100; 
assign wn_re[600] = 26'b11111111111111111011101110; assign wn_im[600] = 26'b11111111111111110000100101; 
assign wn_re[601] = 26'b11111111111111111011101011; assign wn_im[601] = 26'b11111111111111110000100101; 
assign wn_re[602] = 26'b11111111111111111011101000; assign wn_im[602] = 26'b11111111111111110000100110; 
assign wn_re[603] = 26'b11111111111111111011100101; assign wn_im[603] = 26'b11111111111111110000100111; 
assign wn_re[604] = 26'b11111111111111111011100010; assign wn_im[604] = 26'b11111111111111110000101000; 
assign wn_re[605] = 26'b11111111111111111011011111; assign wn_im[605] = 26'b11111111111111110000101001; 
assign wn_re[606] = 26'b11111111111111111011011100; assign wn_im[606] = 26'b11111111111111110000101010; 
assign wn_re[607] = 26'b11111111111111111011011001; assign wn_im[607] = 26'b11111111111111110000101011; 
assign wn_re[608] = 26'b11111111111111111011010110; assign wn_im[608] = 26'b11111111111111110000101100; 
assign wn_re[609] = 26'b11111111111111111011010011; assign wn_im[609] = 26'b11111111111111110000101101; 
assign wn_re[610] = 26'b11111111111111111011010000; assign wn_im[610] = 26'b11111111111111110000101101; 
assign wn_re[611] = 26'b11111111111111111011001101; assign wn_im[611] = 26'b11111111111111110000101110; 
assign wn_re[612] = 26'b11111111111111111011001010; assign wn_im[612] = 26'b11111111111111110000101111; 
assign wn_re[613] = 26'b11111111111111111011000111; assign wn_im[613] = 26'b11111111111111110000110000; 
assign wn_re[614] = 26'b11111111111111111011000100; assign wn_im[614] = 26'b11111111111111110000110001; 
assign wn_re[615] = 26'b11111111111111111011000001; assign wn_im[615] = 26'b11111111111111110000110010; 
assign wn_re[616] = 26'b11111111111111111010111110; assign wn_im[616] = 26'b11111111111111110000110011; 
assign wn_re[617] = 26'b11111111111111111010111011; assign wn_im[617] = 26'b11111111111111110000110100; 
assign wn_re[618] = 26'b11111111111111111010111000; assign wn_im[618] = 26'b11111111111111110000110101; 
assign wn_re[619] = 26'b11111111111111111010110101; assign wn_im[619] = 26'b11111111111111110000110110; 
assign wn_re[620] = 26'b11111111111111111010110010; assign wn_im[620] = 26'b11111111111111110000110111; 
assign wn_re[621] = 26'b11111111111111111010101111; assign wn_im[621] = 26'b11111111111111110000111000; 
assign wn_re[622] = 26'b11111111111111111010101100; assign wn_im[622] = 26'b11111111111111110000111001; 
assign wn_re[623] = 26'b11111111111111111010101001; assign wn_im[623] = 26'b11111111111111110000111010; 
assign wn_re[624] = 26'b11111111111111111010100111; assign wn_im[624] = 26'b11111111111111110000111011; 
assign wn_re[625] = 26'b11111111111111111010100100; assign wn_im[625] = 26'b11111111111111110000111100; 
assign wn_re[626] = 26'b11111111111111111010100001; assign wn_im[626] = 26'b11111111111111110000111101; 
assign wn_re[627] = 26'b11111111111111111010011110; assign wn_im[627] = 26'b11111111111111110000111111; 
assign wn_re[628] = 26'b11111111111111111010011011; assign wn_im[628] = 26'b11111111111111110001000000; 
assign wn_re[629] = 26'b11111111111111111010011000; assign wn_im[629] = 26'b11111111111111110001000001; 
assign wn_re[630] = 26'b11111111111111111010010101; assign wn_im[630] = 26'b11111111111111110001000010; 
assign wn_re[631] = 26'b11111111111111111010010010; assign wn_im[631] = 26'b11111111111111110001000011; 
assign wn_re[632] = 26'b11111111111111111010001111; assign wn_im[632] = 26'b11111111111111110001000100; 
assign wn_re[633] = 26'b11111111111111111010001100; assign wn_im[633] = 26'b11111111111111110001000101; 
assign wn_re[634] = 26'b11111111111111111010001001; assign wn_im[634] = 26'b11111111111111110001000110; 
assign wn_re[635] = 26'b11111111111111111010000110; assign wn_im[635] = 26'b11111111111111110001001000; 
assign wn_re[636] = 26'b11111111111111111010000011; assign wn_im[636] = 26'b11111111111111110001001001; 
assign wn_re[637] = 26'b11111111111111111010000000; assign wn_im[637] = 26'b11111111111111110001001010; 
assign wn_re[638] = 26'b11111111111111111001111101; assign wn_im[638] = 26'b11111111111111110001001011; 
assign wn_re[639] = 26'b11111111111111111001111011; assign wn_im[639] = 26'b11111111111111110001001100; 
assign wn_re[640] = 26'b11111111111111111001111000; assign wn_im[640] = 26'b11111111111111110001001101; 
assign wn_re[641] = 26'b11111111111111111001110101; assign wn_im[641] = 26'b11111111111111110001001111; 
assign wn_re[642] = 26'b11111111111111111001110010; assign wn_im[642] = 26'b11111111111111110001010000; 
assign wn_re[643] = 26'b11111111111111111001101111; assign wn_im[643] = 26'b11111111111111110001010001; 
assign wn_re[644] = 26'b11111111111111111001101100; assign wn_im[644] = 26'b11111111111111110001010010; 
assign wn_re[645] = 26'b11111111111111111001101001; assign wn_im[645] = 26'b11111111111111110001010100; 
assign wn_re[646] = 26'b11111111111111111001100110; assign wn_im[646] = 26'b11111111111111110001010101; 
assign wn_re[647] = 26'b11111111111111111001100011; assign wn_im[647] = 26'b11111111111111110001010110; 
assign wn_re[648] = 26'b11111111111111111001100001; assign wn_im[648] = 26'b11111111111111110001010111; 
assign wn_re[649] = 26'b11111111111111111001011110; assign wn_im[649] = 26'b11111111111111110001011001; 
assign wn_re[650] = 26'b11111111111111111001011011; assign wn_im[650] = 26'b11111111111111110001011010; 
assign wn_re[651] = 26'b11111111111111111001011000; assign wn_im[651] = 26'b11111111111111110001011011; 
assign wn_re[652] = 26'b11111111111111111001010101; assign wn_im[652] = 26'b11111111111111110001011101; 
assign wn_re[653] = 26'b11111111111111111001010010; assign wn_im[653] = 26'b11111111111111110001011110; 
assign wn_re[654] = 26'b11111111111111111001001111; assign wn_im[654] = 26'b11111111111111110001011111; 
assign wn_re[655] = 26'b11111111111111111001001101; assign wn_im[655] = 26'b11111111111111110001100000; 
assign wn_re[656] = 26'b11111111111111111001001010; assign wn_im[656] = 26'b11111111111111110001100010; 
assign wn_re[657] = 26'b11111111111111111001000111; assign wn_im[657] = 26'b11111111111111110001100011; 
assign wn_re[658] = 26'b11111111111111111001000100; assign wn_im[658] = 26'b11111111111111110001100101; 
assign wn_re[659] = 26'b11111111111111111001000001; assign wn_im[659] = 26'b11111111111111110001100110; 
assign wn_re[660] = 26'b11111111111111111000111110; assign wn_im[660] = 26'b11111111111111110001100111; 
assign wn_re[661] = 26'b11111111111111111000111100; assign wn_im[661] = 26'b11111111111111110001101001; 
assign wn_re[662] = 26'b11111111111111111000111001; assign wn_im[662] = 26'b11111111111111110001101010; 
assign wn_re[663] = 26'b11111111111111111000110110; assign wn_im[663] = 26'b11111111111111110001101011; 
assign wn_re[664] = 26'b11111111111111111000110011; assign wn_im[664] = 26'b11111111111111110001101101; 
assign wn_re[665] = 26'b11111111111111111000110000; assign wn_im[665] = 26'b11111111111111110001101110; 
assign wn_re[666] = 26'b11111111111111111000101101; assign wn_im[666] = 26'b11111111111111110001110000; 
assign wn_re[667] = 26'b11111111111111111000101011; assign wn_im[667] = 26'b11111111111111110001110001; 
assign wn_re[668] = 26'b11111111111111111000101000; assign wn_im[668] = 26'b11111111111111110001110011; 
assign wn_re[669] = 26'b11111111111111111000100101; assign wn_im[669] = 26'b11111111111111110001110100; 
assign wn_re[670] = 26'b11111111111111111000100010; assign wn_im[670] = 26'b11111111111111110001110101; 
assign wn_re[671] = 26'b11111111111111111000100000; assign wn_im[671] = 26'b11111111111111110001110111; 
assign wn_re[672] = 26'b11111111111111111000011101; assign wn_im[672] = 26'b11111111111111110001111000; 
assign wn_re[673] = 26'b11111111111111111000011010; assign wn_im[673] = 26'b11111111111111110001111010; 
assign wn_re[674] = 26'b11111111111111111000010111; assign wn_im[674] = 26'b11111111111111110001111011; 
assign wn_re[675] = 26'b11111111111111111000010100; assign wn_im[675] = 26'b11111111111111110001111101; 
assign wn_re[676] = 26'b11111111111111111000010010; assign wn_im[676] = 26'b11111111111111110001111110; 
assign wn_re[677] = 26'b11111111111111111000001111; assign wn_im[677] = 26'b11111111111111110010000000; 
assign wn_re[678] = 26'b11111111111111111000001100; assign wn_im[678] = 26'b11111111111111110010000001; 
assign wn_re[679] = 26'b11111111111111111000001010; assign wn_im[679] = 26'b11111111111111110010000011; 
assign wn_re[680] = 26'b11111111111111111000000111; assign wn_im[680] = 26'b11111111111111110010000101; 
assign wn_re[681] = 26'b11111111111111111000000100; assign wn_im[681] = 26'b11111111111111110010000110; 
assign wn_re[682] = 26'b11111111111111111000000001; assign wn_im[682] = 26'b11111111111111110010001000; 
assign wn_re[683] = 26'b11111111111111110111111111; assign wn_im[683] = 26'b11111111111111110010001001; 
assign wn_re[684] = 26'b11111111111111110111111100; assign wn_im[684] = 26'b11111111111111110010001011; 
assign wn_re[685] = 26'b11111111111111110111111001; assign wn_im[685] = 26'b11111111111111110010001100; 
assign wn_re[686] = 26'b11111111111111110111110110; assign wn_im[686] = 26'b11111111111111110010001110; 
assign wn_re[687] = 26'b11111111111111110111110100; assign wn_im[687] = 26'b11111111111111110010010000; 
assign wn_re[688] = 26'b11111111111111110111110001; assign wn_im[688] = 26'b11111111111111110010010001; 
assign wn_re[689] = 26'b11111111111111110111101110; assign wn_im[689] = 26'b11111111111111110010010011; 
assign wn_re[690] = 26'b11111111111111110111101100; assign wn_im[690] = 26'b11111111111111110010010100; 
assign wn_re[691] = 26'b11111111111111110111101001; assign wn_im[691] = 26'b11111111111111110010010110; 
assign wn_re[692] = 26'b11111111111111110111100110; assign wn_im[692] = 26'b11111111111111110010011000; 
assign wn_re[693] = 26'b11111111111111110111100100; assign wn_im[693] = 26'b11111111111111110010011001; 
assign wn_re[694] = 26'b11111111111111110111100001; assign wn_im[694] = 26'b11111111111111110010011011; 
assign wn_re[695] = 26'b11111111111111110111011110; assign wn_im[695] = 26'b11111111111111110010011101; 
assign wn_re[696] = 26'b11111111111111110111011100; assign wn_im[696] = 26'b11111111111111110010011110; 
assign wn_re[697] = 26'b11111111111111110111011001; assign wn_im[697] = 26'b11111111111111110010100000; 
assign wn_re[698] = 26'b11111111111111110111010110; assign wn_im[698] = 26'b11111111111111110010100010; 
assign wn_re[699] = 26'b11111111111111110111010100; assign wn_im[699] = 26'b11111111111111110010100011; 
assign wn_re[700] = 26'b11111111111111110111010001; assign wn_im[700] = 26'b11111111111111110010100101; 
assign wn_re[701] = 26'b11111111111111110111001110; assign wn_im[701] = 26'b11111111111111110010100111; 
assign wn_re[702] = 26'b11111111111111110111001100; assign wn_im[702] = 26'b11111111111111110010101001; 
assign wn_re[703] = 26'b11111111111111110111001001; assign wn_im[703] = 26'b11111111111111110010101010; 
assign wn_re[704] = 26'b11111111111111110111000111; assign wn_im[704] = 26'b11111111111111110010101100; 
assign wn_re[705] = 26'b11111111111111110111000100; assign wn_im[705] = 26'b11111111111111110010101110; 
assign wn_re[706] = 26'b11111111111111110111000001; assign wn_im[706] = 26'b11111111111111110010110000; 
assign wn_re[707] = 26'b11111111111111110110111111; assign wn_im[707] = 26'b11111111111111110010110001; 
assign wn_re[708] = 26'b11111111111111110110111100; assign wn_im[708] = 26'b11111111111111110010110011; 
assign wn_re[709] = 26'b11111111111111110110111010; assign wn_im[709] = 26'b11111111111111110010110101; 
assign wn_re[710] = 26'b11111111111111110110110111; assign wn_im[710] = 26'b11111111111111110010110111; 
assign wn_re[711] = 26'b11111111111111110110110100; assign wn_im[711] = 26'b11111111111111110010111000; 
assign wn_re[712] = 26'b11111111111111110110110010; assign wn_im[712] = 26'b11111111111111110010111010; 
assign wn_re[713] = 26'b11111111111111110110101111; assign wn_im[713] = 26'b11111111111111110010111100; 
assign wn_re[714] = 26'b11111111111111110110101101; assign wn_im[714] = 26'b11111111111111110010111110; 
assign wn_re[715] = 26'b11111111111111110110101010; assign wn_im[715] = 26'b11111111111111110011000000; 
assign wn_re[716] = 26'b11111111111111110110101000; assign wn_im[716] = 26'b11111111111111110011000010; 
assign wn_re[717] = 26'b11111111111111110110100101; assign wn_im[717] = 26'b11111111111111110011000011; 
assign wn_re[718] = 26'b11111111111111110110100011; assign wn_im[718] = 26'b11111111111111110011000101; 
assign wn_re[719] = 26'b11111111111111110110100000; assign wn_im[719] = 26'b11111111111111110011000111; 
assign wn_re[720] = 26'b11111111111111110110011110; assign wn_im[720] = 26'b11111111111111110011001001; 
assign wn_re[721] = 26'b11111111111111110110011011; assign wn_im[721] = 26'b11111111111111110011001011; 
assign wn_re[722] = 26'b11111111111111110110011000; assign wn_im[722] = 26'b11111111111111110011001101; 
assign wn_re[723] = 26'b11111111111111110110010110; assign wn_im[723] = 26'b11111111111111110011001111; 
assign wn_re[724] = 26'b11111111111111110110010011; assign wn_im[724] = 26'b11111111111111110011010001; 
assign wn_re[725] = 26'b11111111111111110110010001; assign wn_im[725] = 26'b11111111111111110011010010; 
assign wn_re[726] = 26'b11111111111111110110001110; assign wn_im[726] = 26'b11111111111111110011010100; 
assign wn_re[727] = 26'b11111111111111110110001100; assign wn_im[727] = 26'b11111111111111110011010110; 
assign wn_re[728] = 26'b11111111111111110110001010; assign wn_im[728] = 26'b11111111111111110011011000; 
assign wn_re[729] = 26'b11111111111111110110000111; assign wn_im[729] = 26'b11111111111111110011011010; 
assign wn_re[730] = 26'b11111111111111110110000101; assign wn_im[730] = 26'b11111111111111110011011100; 
assign wn_re[731] = 26'b11111111111111110110000010; assign wn_im[731] = 26'b11111111111111110011011110; 
assign wn_re[732] = 26'b11111111111111110110000000; assign wn_im[732] = 26'b11111111111111110011100000; 
assign wn_re[733] = 26'b11111111111111110101111101; assign wn_im[733] = 26'b11111111111111110011100010; 
assign wn_re[734] = 26'b11111111111111110101111011; assign wn_im[734] = 26'b11111111111111110011100100; 
assign wn_re[735] = 26'b11111111111111110101111000; assign wn_im[735] = 26'b11111111111111110011100110; 
assign wn_re[736] = 26'b11111111111111110101110110; assign wn_im[736] = 26'b11111111111111110011101000; 
assign wn_re[737] = 26'b11111111111111110101110011; assign wn_im[737] = 26'b11111111111111110011101010; 
assign wn_re[738] = 26'b11111111111111110101110001; assign wn_im[738] = 26'b11111111111111110011101100; 
assign wn_re[739] = 26'b11111111111111110101101111; assign wn_im[739] = 26'b11111111111111110011101110; 
assign wn_re[740] = 26'b11111111111111110101101100; assign wn_im[740] = 26'b11111111111111110011110000; 
assign wn_re[741] = 26'b11111111111111110101101010; assign wn_im[741] = 26'b11111111111111110011110010; 
assign wn_re[742] = 26'b11111111111111110101100111; assign wn_im[742] = 26'b11111111111111110011110100; 
assign wn_re[743] = 26'b11111111111111110101100101; assign wn_im[743] = 26'b11111111111111110011110110; 
assign wn_re[744] = 26'b11111111111111110101100011; assign wn_im[744] = 26'b11111111111111110011111000; 
assign wn_re[745] = 26'b11111111111111110101100000; assign wn_im[745] = 26'b11111111111111110011111010; 
assign wn_re[746] = 26'b11111111111111110101011110; assign wn_im[746] = 26'b11111111111111110011111100; 
assign wn_re[747] = 26'b11111111111111110101011100; assign wn_im[747] = 26'b11111111111111110011111110; 
assign wn_re[748] = 26'b11111111111111110101011001; assign wn_im[748] = 26'b11111111111111110100000000; 
assign wn_re[749] = 26'b11111111111111110101010111; assign wn_im[749] = 26'b11111111111111110100000010; 
assign wn_re[750] = 26'b11111111111111110101010100; assign wn_im[750] = 26'b11111111111111110100000101; 
assign wn_re[751] = 26'b11111111111111110101010010; assign wn_im[751] = 26'b11111111111111110100000111; 
assign wn_re[752] = 26'b11111111111111110101010000; assign wn_im[752] = 26'b11111111111111110100001001; 
assign wn_re[753] = 26'b11111111111111110101001101; assign wn_im[753] = 26'b11111111111111110100001011; 
assign wn_re[754] = 26'b11111111111111110101001011; assign wn_im[754] = 26'b11111111111111110100001101; 
assign wn_re[755] = 26'b11111111111111110101001001; assign wn_im[755] = 26'b11111111111111110100001111; 
assign wn_re[756] = 26'b11111111111111110101000111; assign wn_im[756] = 26'b11111111111111110100010001; 
assign wn_re[757] = 26'b11111111111111110101000100; assign wn_im[757] = 26'b11111111111111110100010011; 
assign wn_re[758] = 26'b11111111111111110101000010; assign wn_im[758] = 26'b11111111111111110100010110; 
assign wn_re[759] = 26'b11111111111111110101000000; assign wn_im[759] = 26'b11111111111111110100011000; 
assign wn_re[760] = 26'b11111111111111110100111101; assign wn_im[760] = 26'b11111111111111110100011010; 
assign wn_re[761] = 26'b11111111111111110100111011; assign wn_im[761] = 26'b11111111111111110100011100; 
assign wn_re[762] = 26'b11111111111111110100111001; assign wn_im[762] = 26'b11111111111111110100011110; 
assign wn_re[763] = 26'b11111111111111110100110111; assign wn_im[763] = 26'b11111111111111110100100000; 
assign wn_re[764] = 26'b11111111111111110100110100; assign wn_im[764] = 26'b11111111111111110100100011; 
assign wn_re[765] = 26'b11111111111111110100110010; assign wn_im[765] = 26'b11111111111111110100100101; 
assign wn_re[766] = 26'b11111111111111110100110000; assign wn_im[766] = 26'b11111111111111110100100111; 
assign wn_re[767] = 26'b11111111111111110100101110; assign wn_im[767] = 26'b11111111111111110100101001; 
assign wn_re[768] = 26'b11111111111111110100101011; assign wn_im[768] = 26'b11111111111111110100101011; 
assign wn_re[769] = 26'b11111111111111110100101001; assign wn_im[769] = 26'b11111111111111110100101110; 
assign wn_re[770] = 26'b11111111111111110100100111; assign wn_im[770] = 26'b11111111111111110100110000; 
assign wn_re[771] = 26'b11111111111111110100100101; assign wn_im[771] = 26'b11111111111111110100110010; 
assign wn_re[772] = 26'b11111111111111110100100011; assign wn_im[772] = 26'b11111111111111110100110100; 
assign wn_re[773] = 26'b11111111111111110100100000; assign wn_im[773] = 26'b11111111111111110100110111; 
assign wn_re[774] = 26'b11111111111111110100011110; assign wn_im[774] = 26'b11111111111111110100111001; 
assign wn_re[775] = 26'b11111111111111110100011100; assign wn_im[775] = 26'b11111111111111110100111011; 
assign wn_re[776] = 26'b11111111111111110100011010; assign wn_im[776] = 26'b11111111111111110100111101; 
assign wn_re[777] = 26'b11111111111111110100011000; assign wn_im[777] = 26'b11111111111111110101000000; 
assign wn_re[778] = 26'b11111111111111110100010110; assign wn_im[778] = 26'b11111111111111110101000010; 
assign wn_re[779] = 26'b11111111111111110100010011; assign wn_im[779] = 26'b11111111111111110101000100; 
assign wn_re[780] = 26'b11111111111111110100010001; assign wn_im[780] = 26'b11111111111111110101000111; 
assign wn_re[781] = 26'b11111111111111110100001111; assign wn_im[781] = 26'b11111111111111110101001001; 
assign wn_re[782] = 26'b11111111111111110100001101; assign wn_im[782] = 26'b11111111111111110101001011; 
assign wn_re[783] = 26'b11111111111111110100001011; assign wn_im[783] = 26'b11111111111111110101001101; 
assign wn_re[784] = 26'b11111111111111110100001001; assign wn_im[784] = 26'b11111111111111110101010000; 
assign wn_re[785] = 26'b11111111111111110100000111; assign wn_im[785] = 26'b11111111111111110101010010; 
assign wn_re[786] = 26'b11111111111111110100000101; assign wn_im[786] = 26'b11111111111111110101010100; 
assign wn_re[787] = 26'b11111111111111110100000010; assign wn_im[787] = 26'b11111111111111110101010111; 
assign wn_re[788] = 26'b11111111111111110100000000; assign wn_im[788] = 26'b11111111111111110101011001; 
assign wn_re[789] = 26'b11111111111111110011111110; assign wn_im[789] = 26'b11111111111111110101011100; 
assign wn_re[790] = 26'b11111111111111110011111100; assign wn_im[790] = 26'b11111111111111110101011110; 
assign wn_re[791] = 26'b11111111111111110011111010; assign wn_im[791] = 26'b11111111111111110101100000; 
assign wn_re[792] = 26'b11111111111111110011111000; assign wn_im[792] = 26'b11111111111111110101100011; 
assign wn_re[793] = 26'b11111111111111110011110110; assign wn_im[793] = 26'b11111111111111110101100101; 
assign wn_re[794] = 26'b11111111111111110011110100; assign wn_im[794] = 26'b11111111111111110101100111; 
assign wn_re[795] = 26'b11111111111111110011110010; assign wn_im[795] = 26'b11111111111111110101101010; 
assign wn_re[796] = 26'b11111111111111110011110000; assign wn_im[796] = 26'b11111111111111110101101100; 
assign wn_re[797] = 26'b11111111111111110011101110; assign wn_im[797] = 26'b11111111111111110101101111; 
assign wn_re[798] = 26'b11111111111111110011101100; assign wn_im[798] = 26'b11111111111111110101110001; 
assign wn_re[799] = 26'b11111111111111110011101010; assign wn_im[799] = 26'b11111111111111110101110011; 
assign wn_re[800] = 26'b11111111111111110011101000; assign wn_im[800] = 26'b11111111111111110101110110; 
assign wn_re[801] = 26'b11111111111111110011100110; assign wn_im[801] = 26'b11111111111111110101111000; 
assign wn_re[802] = 26'b11111111111111110011100100; assign wn_im[802] = 26'b11111111111111110101111011; 
assign wn_re[803] = 26'b11111111111111110011100010; assign wn_im[803] = 26'b11111111111111110101111101; 
assign wn_re[804] = 26'b11111111111111110011100000; assign wn_im[804] = 26'b11111111111111110110000000; 
assign wn_re[805] = 26'b11111111111111110011011110; assign wn_im[805] = 26'b11111111111111110110000010; 
assign wn_re[806] = 26'b11111111111111110011011100; assign wn_im[806] = 26'b11111111111111110110000101; 
assign wn_re[807] = 26'b11111111111111110011011010; assign wn_im[807] = 26'b11111111111111110110000111; 
assign wn_re[808] = 26'b11111111111111110011011000; assign wn_im[808] = 26'b11111111111111110110001010; 
assign wn_re[809] = 26'b11111111111111110011010110; assign wn_im[809] = 26'b11111111111111110110001100; 
assign wn_re[810] = 26'b11111111111111110011010100; assign wn_im[810] = 26'b11111111111111110110001110; 
assign wn_re[811] = 26'b11111111111111110011010010; assign wn_im[811] = 26'b11111111111111110110010001; 
assign wn_re[812] = 26'b11111111111111110011010001; assign wn_im[812] = 26'b11111111111111110110010011; 
assign wn_re[813] = 26'b11111111111111110011001111; assign wn_im[813] = 26'b11111111111111110110010110; 
assign wn_re[814] = 26'b11111111111111110011001101; assign wn_im[814] = 26'b11111111111111110110011000; 
assign wn_re[815] = 26'b11111111111111110011001011; assign wn_im[815] = 26'b11111111111111110110011011; 
assign wn_re[816] = 26'b11111111111111110011001001; assign wn_im[816] = 26'b11111111111111110110011110; 
assign wn_re[817] = 26'b11111111111111110011000111; assign wn_im[817] = 26'b11111111111111110110100000; 
assign wn_re[818] = 26'b11111111111111110011000101; assign wn_im[818] = 26'b11111111111111110110100011; 
assign wn_re[819] = 26'b11111111111111110011000011; assign wn_im[819] = 26'b11111111111111110110100101; 
assign wn_re[820] = 26'b11111111111111110011000010; assign wn_im[820] = 26'b11111111111111110110101000; 
assign wn_re[821] = 26'b11111111111111110011000000; assign wn_im[821] = 26'b11111111111111110110101010; 
assign wn_re[822] = 26'b11111111111111110010111110; assign wn_im[822] = 26'b11111111111111110110101101; 
assign wn_re[823] = 26'b11111111111111110010111100; assign wn_im[823] = 26'b11111111111111110110101111; 
assign wn_re[824] = 26'b11111111111111110010111010; assign wn_im[824] = 26'b11111111111111110110110010; 
assign wn_re[825] = 26'b11111111111111110010111000; assign wn_im[825] = 26'b11111111111111110110110100; 
assign wn_re[826] = 26'b11111111111111110010110111; assign wn_im[826] = 26'b11111111111111110110110111; 
assign wn_re[827] = 26'b11111111111111110010110101; assign wn_im[827] = 26'b11111111111111110110111010; 
assign wn_re[828] = 26'b11111111111111110010110011; assign wn_im[828] = 26'b11111111111111110110111100; 
assign wn_re[829] = 26'b11111111111111110010110001; assign wn_im[829] = 26'b11111111111111110110111111; 
assign wn_re[830] = 26'b11111111111111110010110000; assign wn_im[830] = 26'b11111111111111110111000001; 
assign wn_re[831] = 26'b11111111111111110010101110; assign wn_im[831] = 26'b11111111111111110111000100; 
assign wn_re[832] = 26'b11111111111111110010101100; assign wn_im[832] = 26'b11111111111111110111000111; 
assign wn_re[833] = 26'b11111111111111110010101010; assign wn_im[833] = 26'b11111111111111110111001001; 
assign wn_re[834] = 26'b11111111111111110010101001; assign wn_im[834] = 26'b11111111111111110111001100; 
assign wn_re[835] = 26'b11111111111111110010100111; assign wn_im[835] = 26'b11111111111111110111001110; 
assign wn_re[836] = 26'b11111111111111110010100101; assign wn_im[836] = 26'b11111111111111110111010001; 
assign wn_re[837] = 26'b11111111111111110010100011; assign wn_im[837] = 26'b11111111111111110111010100; 
assign wn_re[838] = 26'b11111111111111110010100010; assign wn_im[838] = 26'b11111111111111110111010110; 
assign wn_re[839] = 26'b11111111111111110010100000; assign wn_im[839] = 26'b11111111111111110111011001; 
assign wn_re[840] = 26'b11111111111111110010011110; assign wn_im[840] = 26'b11111111111111110111011100; 
assign wn_re[841] = 26'b11111111111111110010011101; assign wn_im[841] = 26'b11111111111111110111011110; 
assign wn_re[842] = 26'b11111111111111110010011011; assign wn_im[842] = 26'b11111111111111110111100001; 
assign wn_re[843] = 26'b11111111111111110010011001; assign wn_im[843] = 26'b11111111111111110111100100; 
assign wn_re[844] = 26'b11111111111111110010011000; assign wn_im[844] = 26'b11111111111111110111100110; 
assign wn_re[845] = 26'b11111111111111110010010110; assign wn_im[845] = 26'b11111111111111110111101001; 
assign wn_re[846] = 26'b11111111111111110010010100; assign wn_im[846] = 26'b11111111111111110111101100; 
assign wn_re[847] = 26'b11111111111111110010010011; assign wn_im[847] = 26'b11111111111111110111101110; 
assign wn_re[848] = 26'b11111111111111110010010001; assign wn_im[848] = 26'b11111111111111110111110001; 
assign wn_re[849] = 26'b11111111111111110010010000; assign wn_im[849] = 26'b11111111111111110111110100; 
assign wn_re[850] = 26'b11111111111111110010001110; assign wn_im[850] = 26'b11111111111111110111110110; 
assign wn_re[851] = 26'b11111111111111110010001100; assign wn_im[851] = 26'b11111111111111110111111001; 
assign wn_re[852] = 26'b11111111111111110010001011; assign wn_im[852] = 26'b11111111111111110111111100; 
assign wn_re[853] = 26'b11111111111111110010001001; assign wn_im[853] = 26'b11111111111111110111111111; 
assign wn_re[854] = 26'b11111111111111110010001000; assign wn_im[854] = 26'b11111111111111111000000001; 
assign wn_re[855] = 26'b11111111111111110010000110; assign wn_im[855] = 26'b11111111111111111000000100; 
assign wn_re[856] = 26'b11111111111111110010000101; assign wn_im[856] = 26'b11111111111111111000000111; 
assign wn_re[857] = 26'b11111111111111110010000011; assign wn_im[857] = 26'b11111111111111111000001010; 
assign wn_re[858] = 26'b11111111111111110010000001; assign wn_im[858] = 26'b11111111111111111000001100; 
assign wn_re[859] = 26'b11111111111111110010000000; assign wn_im[859] = 26'b11111111111111111000001111; 
assign wn_re[860] = 26'b11111111111111110001111110; assign wn_im[860] = 26'b11111111111111111000010010; 
assign wn_re[861] = 26'b11111111111111110001111101; assign wn_im[861] = 26'b11111111111111111000010100; 
assign wn_re[862] = 26'b11111111111111110001111011; assign wn_im[862] = 26'b11111111111111111000010111; 
assign wn_re[863] = 26'b11111111111111110001111010; assign wn_im[863] = 26'b11111111111111111000011010; 
assign wn_re[864] = 26'b11111111111111110001111000; assign wn_im[864] = 26'b11111111111111111000011101; 
assign wn_re[865] = 26'b11111111111111110001110111; assign wn_im[865] = 26'b11111111111111111000100000; 
assign wn_re[866] = 26'b11111111111111110001110101; assign wn_im[866] = 26'b11111111111111111000100010; 
assign wn_re[867] = 26'b11111111111111110001110100; assign wn_im[867] = 26'b11111111111111111000100101; 
assign wn_re[868] = 26'b11111111111111110001110011; assign wn_im[868] = 26'b11111111111111111000101000; 
assign wn_re[869] = 26'b11111111111111110001110001; assign wn_im[869] = 26'b11111111111111111000101011; 
assign wn_re[870] = 26'b11111111111111110001110000; assign wn_im[870] = 26'b11111111111111111000101101; 
assign wn_re[871] = 26'b11111111111111110001101110; assign wn_im[871] = 26'b11111111111111111000110000; 
assign wn_re[872] = 26'b11111111111111110001101101; assign wn_im[872] = 26'b11111111111111111000110011; 
assign wn_re[873] = 26'b11111111111111110001101011; assign wn_im[873] = 26'b11111111111111111000110110; 
assign wn_re[874] = 26'b11111111111111110001101010; assign wn_im[874] = 26'b11111111111111111000111001; 
assign wn_re[875] = 26'b11111111111111110001101001; assign wn_im[875] = 26'b11111111111111111000111100; 
assign wn_re[876] = 26'b11111111111111110001100111; assign wn_im[876] = 26'b11111111111111111000111110; 
assign wn_re[877] = 26'b11111111111111110001100110; assign wn_im[877] = 26'b11111111111111111001000001; 
assign wn_re[878] = 26'b11111111111111110001100101; assign wn_im[878] = 26'b11111111111111111001000100; 
assign wn_re[879] = 26'b11111111111111110001100011; assign wn_im[879] = 26'b11111111111111111001000111; 
assign wn_re[880] = 26'b11111111111111110001100010; assign wn_im[880] = 26'b11111111111111111001001010; 
assign wn_re[881] = 26'b11111111111111110001100000; assign wn_im[881] = 26'b11111111111111111001001101; 
assign wn_re[882] = 26'b11111111111111110001011111; assign wn_im[882] = 26'b11111111111111111001001111; 
assign wn_re[883] = 26'b11111111111111110001011110; assign wn_im[883] = 26'b11111111111111111001010010; 
assign wn_re[884] = 26'b11111111111111110001011101; assign wn_im[884] = 26'b11111111111111111001010101; 
assign wn_re[885] = 26'b11111111111111110001011011; assign wn_im[885] = 26'b11111111111111111001011000; 
assign wn_re[886] = 26'b11111111111111110001011010; assign wn_im[886] = 26'b11111111111111111001011011; 
assign wn_re[887] = 26'b11111111111111110001011001; assign wn_im[887] = 26'b11111111111111111001011110; 
assign wn_re[888] = 26'b11111111111111110001010111; assign wn_im[888] = 26'b11111111111111111001100001; 
assign wn_re[889] = 26'b11111111111111110001010110; assign wn_im[889] = 26'b11111111111111111001100011; 
assign wn_re[890] = 26'b11111111111111110001010101; assign wn_im[890] = 26'b11111111111111111001100110; 
assign wn_re[891] = 26'b11111111111111110001010100; assign wn_im[891] = 26'b11111111111111111001101001; 
assign wn_re[892] = 26'b11111111111111110001010010; assign wn_im[892] = 26'b11111111111111111001101100; 
assign wn_re[893] = 26'b11111111111111110001010001; assign wn_im[893] = 26'b11111111111111111001101111; 
assign wn_re[894] = 26'b11111111111111110001010000; assign wn_im[894] = 26'b11111111111111111001110010; 
assign wn_re[895] = 26'b11111111111111110001001111; assign wn_im[895] = 26'b11111111111111111001110101; 
assign wn_re[896] = 26'b11111111111111110001001101; assign wn_im[896] = 26'b11111111111111111001111000; 
assign wn_re[897] = 26'b11111111111111110001001100; assign wn_im[897] = 26'b11111111111111111001111011; 
assign wn_re[898] = 26'b11111111111111110001001011; assign wn_im[898] = 26'b11111111111111111001111101; 
assign wn_re[899] = 26'b11111111111111110001001010; assign wn_im[899] = 26'b11111111111111111010000000; 
assign wn_re[900] = 26'b11111111111111110001001001; assign wn_im[900] = 26'b11111111111111111010000011; 
assign wn_re[901] = 26'b11111111111111110001001000; assign wn_im[901] = 26'b11111111111111111010000110; 
assign wn_re[902] = 26'b11111111111111110001000110; assign wn_im[902] = 26'b11111111111111111010001001; 
assign wn_re[903] = 26'b11111111111111110001000101; assign wn_im[903] = 26'b11111111111111111010001100; 
assign wn_re[904] = 26'b11111111111111110001000100; assign wn_im[904] = 26'b11111111111111111010001111; 
assign wn_re[905] = 26'b11111111111111110001000011; assign wn_im[905] = 26'b11111111111111111010010010; 
assign wn_re[906] = 26'b11111111111111110001000010; assign wn_im[906] = 26'b11111111111111111010010101; 
assign wn_re[907] = 26'b11111111111111110001000001; assign wn_im[907] = 26'b11111111111111111010011000; 
assign wn_re[908] = 26'b11111111111111110001000000; assign wn_im[908] = 26'b11111111111111111010011011; 
assign wn_re[909] = 26'b11111111111111110000111111; assign wn_im[909] = 26'b11111111111111111010011110; 
assign wn_re[910] = 26'b11111111111111110000111101; assign wn_im[910] = 26'b11111111111111111010100001; 
assign wn_re[911] = 26'b11111111111111110000111100; assign wn_im[911] = 26'b11111111111111111010100100; 
assign wn_re[912] = 26'b11111111111111110000111011; assign wn_im[912] = 26'b11111111111111111010100111; 
assign wn_re[913] = 26'b11111111111111110000111010; assign wn_im[913] = 26'b11111111111111111010101001; 
assign wn_re[914] = 26'b11111111111111110000111001; assign wn_im[914] = 26'b11111111111111111010101100; 
assign wn_re[915] = 26'b11111111111111110000111000; assign wn_im[915] = 26'b11111111111111111010101111; 
assign wn_re[916] = 26'b11111111111111110000110111; assign wn_im[916] = 26'b11111111111111111010110010; 
assign wn_re[917] = 26'b11111111111111110000110110; assign wn_im[917] = 26'b11111111111111111010110101; 
assign wn_re[918] = 26'b11111111111111110000110101; assign wn_im[918] = 26'b11111111111111111010111000; 
assign wn_re[919] = 26'b11111111111111110000110100; assign wn_im[919] = 26'b11111111111111111010111011; 
assign wn_re[920] = 26'b11111111111111110000110011; assign wn_im[920] = 26'b11111111111111111010111110; 
assign wn_re[921] = 26'b11111111111111110000110010; assign wn_im[921] = 26'b11111111111111111011000001; 
assign wn_re[922] = 26'b11111111111111110000110001; assign wn_im[922] = 26'b11111111111111111011000100; 
assign wn_re[923] = 26'b11111111111111110000110000; assign wn_im[923] = 26'b11111111111111111011000111; 
assign wn_re[924] = 26'b11111111111111110000101111; assign wn_im[924] = 26'b11111111111111111011001010; 
assign wn_re[925] = 26'b11111111111111110000101110; assign wn_im[925] = 26'b11111111111111111011001101; 
assign wn_re[926] = 26'b11111111111111110000101101; assign wn_im[926] = 26'b11111111111111111011010000; 
assign wn_re[927] = 26'b11111111111111110000101101; assign wn_im[927] = 26'b11111111111111111011010011; 
assign wn_re[928] = 26'b11111111111111110000101100; assign wn_im[928] = 26'b11111111111111111011010110; 
assign wn_re[929] = 26'b11111111111111110000101011; assign wn_im[929] = 26'b11111111111111111011011001; 
assign wn_re[930] = 26'b11111111111111110000101010; assign wn_im[930] = 26'b11111111111111111011011100; 
assign wn_re[931] = 26'b11111111111111110000101001; assign wn_im[931] = 26'b11111111111111111011011111; 
assign wn_re[932] = 26'b11111111111111110000101000; assign wn_im[932] = 26'b11111111111111111011100010; 
assign wn_re[933] = 26'b11111111111111110000100111; assign wn_im[933] = 26'b11111111111111111011100101; 
assign wn_re[934] = 26'b11111111111111110000100110; assign wn_im[934] = 26'b11111111111111111011101000; 
assign wn_re[935] = 26'b11111111111111110000100101; assign wn_im[935] = 26'b11111111111111111011101011; 
assign wn_re[936] = 26'b11111111111111110000100101; assign wn_im[936] = 26'b11111111111111111011101110; 
assign wn_re[937] = 26'b11111111111111110000100100; assign wn_im[937] = 26'b11111111111111111011110001; 
assign wn_re[938] = 26'b11111111111111110000100011; assign wn_im[938] = 26'b11111111111111111011110100; 
assign wn_re[939] = 26'b11111111111111110000100010; assign wn_im[939] = 26'b11111111111111111011110111; 
assign wn_re[940] = 26'b11111111111111110000100001; assign wn_im[940] = 26'b11111111111111111011111011; 
assign wn_re[941] = 26'b11111111111111110000100001; assign wn_im[941] = 26'b11111111111111111011111110; 
assign wn_re[942] = 26'b11111111111111110000100000; assign wn_im[942] = 26'b11111111111111111100000001; 
assign wn_re[943] = 26'b11111111111111110000011111; assign wn_im[943] = 26'b11111111111111111100000100; 
assign wn_re[944] = 26'b11111111111111110000011110; assign wn_im[944] = 26'b11111111111111111100000111; 
assign wn_re[945] = 26'b11111111111111110000011101; assign wn_im[945] = 26'b11111111111111111100001010; 
assign wn_re[946] = 26'b11111111111111110000011101; assign wn_im[946] = 26'b11111111111111111100001101; 
assign wn_re[947] = 26'b11111111111111110000011100; assign wn_im[947] = 26'b11111111111111111100010000; 
assign wn_re[948] = 26'b11111111111111110000011011; assign wn_im[948] = 26'b11111111111111111100010011; 
assign wn_re[949] = 26'b11111111111111110000011010; assign wn_im[949] = 26'b11111111111111111100010110; 
assign wn_re[950] = 26'b11111111111111110000011010; assign wn_im[950] = 26'b11111111111111111100011001; 
assign wn_re[951] = 26'b11111111111111110000011001; assign wn_im[951] = 26'b11111111111111111100011100; 
assign wn_re[952] = 26'b11111111111111110000011000; assign wn_im[952] = 26'b11111111111111111100011111; 
assign wn_re[953] = 26'b11111111111111110000011000; assign wn_im[953] = 26'b11111111111111111100100010; 
assign wn_re[954] = 26'b11111111111111110000010111; assign wn_im[954] = 26'b11111111111111111100100101; 
assign wn_re[955] = 26'b11111111111111110000010110; assign wn_im[955] = 26'b11111111111111111100101000; 
assign wn_re[956] = 26'b11111111111111110000010110; assign wn_im[956] = 26'b11111111111111111100101011; 
assign wn_re[957] = 26'b11111111111111110000010101; assign wn_im[957] = 26'b11111111111111111100101110; 
assign wn_re[958] = 26'b11111111111111110000010100; assign wn_im[958] = 26'b11111111111111111100110010; 
assign wn_re[959] = 26'b11111111111111110000010100; assign wn_im[959] = 26'b11111111111111111100110101; 
assign wn_re[960] = 26'b11111111111111110000010011; assign wn_im[960] = 26'b11111111111111111100111000; 
assign wn_re[961] = 26'b11111111111111110000010011; assign wn_im[961] = 26'b11111111111111111100111011; 
assign wn_re[962] = 26'b11111111111111110000010010; assign wn_im[962] = 26'b11111111111111111100111110; 
assign wn_re[963] = 26'b11111111111111110000010001; assign wn_im[963] = 26'b11111111111111111101000001; 
assign wn_re[964] = 26'b11111111111111110000010001; assign wn_im[964] = 26'b11111111111111111101000100; 
assign wn_re[965] = 26'b11111111111111110000010000; assign wn_im[965] = 26'b11111111111111111101000111; 
assign wn_re[966] = 26'b11111111111111110000010000; assign wn_im[966] = 26'b11111111111111111101001010; 
assign wn_re[967] = 26'b11111111111111110000001111; assign wn_im[967] = 26'b11111111111111111101001101; 
assign wn_re[968] = 26'b11111111111111110000001111; assign wn_im[968] = 26'b11111111111111111101010000; 
assign wn_re[969] = 26'b11111111111111110000001110; assign wn_im[969] = 26'b11111111111111111101010100; 
assign wn_re[970] = 26'b11111111111111110000001110; assign wn_im[970] = 26'b11111111111111111101010111; 
assign wn_re[971] = 26'b11111111111111110000001101; assign wn_im[971] = 26'b11111111111111111101011010; 
assign wn_re[972] = 26'b11111111111111110000001101; assign wn_im[972] = 26'b11111111111111111101011101; 
assign wn_re[973] = 26'b11111111111111110000001100; assign wn_im[973] = 26'b11111111111111111101100000; 
assign wn_re[974] = 26'b11111111111111110000001100; assign wn_im[974] = 26'b11111111111111111101100011; 
assign wn_re[975] = 26'b11111111111111110000001011; assign wn_im[975] = 26'b11111111111111111101100110; 
assign wn_re[976] = 26'b11111111111111110000001011; assign wn_im[976] = 26'b11111111111111111101101001; 
assign wn_re[977] = 26'b11111111111111110000001010; assign wn_im[977] = 26'b11111111111111111101101100; 
assign wn_re[978] = 26'b11111111111111110000001010; assign wn_im[978] = 26'b11111111111111111101101111; 
assign wn_re[979] = 26'b11111111111111110000001001; assign wn_im[979] = 26'b11111111111111111101110011; 
assign wn_re[980] = 26'b11111111111111110000001001; assign wn_im[980] = 26'b11111111111111111101110110; 
assign wn_re[981] = 26'b11111111111111110000001000; assign wn_im[981] = 26'b11111111111111111101111001; 
assign wn_re[982] = 26'b11111111111111110000001000; assign wn_im[982] = 26'b11111111111111111101111100; 
assign wn_re[983] = 26'b11111111111111110000001000; assign wn_im[983] = 26'b11111111111111111101111111; 
assign wn_re[984] = 26'b11111111111111110000000111; assign wn_im[984] = 26'b11111111111111111110000010; 
assign wn_re[985] = 26'b11111111111111110000000111; assign wn_im[985] = 26'b11111111111111111110000101; 
assign wn_re[986] = 26'b11111111111111110000000110; assign wn_im[986] = 26'b11111111111111111110001000; 
assign wn_re[987] = 26'b11111111111111110000000110; assign wn_im[987] = 26'b11111111111111111110001100; 
assign wn_re[988] = 26'b11111111111111110000000110; assign wn_im[988] = 26'b11111111111111111110001111; 
assign wn_re[989] = 26'b11111111111111110000000101; assign wn_im[989] = 26'b11111111111111111110010010; 
assign wn_re[990] = 26'b11111111111111110000000101; assign wn_im[990] = 26'b11111111111111111110010101; 
assign wn_re[991] = 26'b11111111111111110000000101; assign wn_im[991] = 26'b11111111111111111110011000; 
assign wn_re[992] = 26'b11111111111111110000000100; assign wn_im[992] = 26'b11111111111111111110011011; 
assign wn_re[993] = 26'b11111111111111110000000100; assign wn_im[993] = 26'b11111111111111111110011110; 
assign wn_re[994] = 26'b11111111111111110000000100; assign wn_im[994] = 26'b11111111111111111110100001; 
assign wn_re[995] = 26'b11111111111111110000000100; assign wn_im[995] = 26'b11111111111111111110100101; 
assign wn_re[996] = 26'b11111111111111110000000011; assign wn_im[996] = 26'b11111111111111111110101000; 
assign wn_re[997] = 26'b11111111111111110000000011; assign wn_im[997] = 26'b11111111111111111110101011; 
assign wn_re[998] = 26'b11111111111111110000000011; assign wn_im[998] = 26'b11111111111111111110101110; 
assign wn_re[999] = 26'b11111111111111110000000011; assign wn_im[999] = 26'b11111111111111111110110001; 
assign wn_re[1000] = 26'b11111111111111110000000010; assign wn_im[1000] = 26'b11111111111111111110110100; 
assign wn_re[1001] = 26'b11111111111111110000000010; assign wn_im[1001] = 26'b11111111111111111110110111; 
assign wn_re[1002] = 26'b11111111111111110000000010; assign wn_im[1002] = 26'b11111111111111111110111010; 
assign wn_re[1003] = 26'b11111111111111110000000010; assign wn_im[1003] = 26'b11111111111111111110111110; 
assign wn_re[1004] = 26'b11111111111111110000000001; assign wn_im[1004] = 26'b11111111111111111111000001; 
assign wn_re[1005] = 26'b11111111111111110000000001; assign wn_im[1005] = 26'b11111111111111111111000100; 
assign wn_re[1006] = 26'b11111111111111110000000001; assign wn_im[1006] = 26'b11111111111111111111000111; 
assign wn_re[1007] = 26'b11111111111111110000000001; assign wn_im[1007] = 26'b11111111111111111111001010; 
assign wn_re[1008] = 26'b11111111111111110000000001; assign wn_im[1008] = 26'b11111111111111111111001101; 
assign wn_re[1009] = 26'b11111111111111110000000001; assign wn_im[1009] = 26'b11111111111111111111010000; 
assign wn_re[1010] = 26'b11111111111111110000000000; assign wn_im[1010] = 26'b11111111111111111111010100; 
assign wn_re[1011] = 26'b11111111111111110000000000; assign wn_im[1011] = 26'b11111111111111111111010111; 
assign wn_re[1012] = 26'b11111111111111110000000000; assign wn_im[1012] = 26'b11111111111111111111011010; 
assign wn_re[1013] = 26'b11111111111111110000000000; assign wn_im[1013] = 26'b11111111111111111111011101; 
assign wn_re[1014] = 26'b11111111111111110000000000; assign wn_im[1014] = 26'b11111111111111111111100000; 
assign wn_re[1015] = 26'b11111111111111110000000000; assign wn_im[1015] = 26'b11111111111111111111100011; 
assign wn_re[1016] = 26'b11111111111111110000000000; assign wn_im[1016] = 26'b11111111111111111111100110; 
assign wn_re[1017] = 26'b11111111111111110000000000; assign wn_im[1017] = 26'b11111111111111111111101010; 
assign wn_re[1018] = 26'b11111111111111110000000000; assign wn_im[1018] = 26'b11111111111111111111101101; 
assign wn_re[1019] = 26'b11111111111111110000000000; assign wn_im[1019] = 26'b11111111111111111111110000; 
assign wn_re[1020] = 26'b11111111111111110000000000; assign wn_im[1020] = 26'b11111111111111111111110011; 
assign wn_re[1021] = 26'b11111111111111110000000000; assign wn_im[1021] = 26'b11111111111111111111110110; 
assign wn_re[1022] = 26'b11111111111111110000000000; assign wn_im[1022] = 26'b11111111111111111111111001; 
assign wn_re[1023] = 26'b11111111111111110000000000; assign wn_im[1023] = 26'b11111111111111111111111100; 
assign wn_re[1024] = 26'b11111111111111110000000000; assign wn_im[1024] = 26'b11111111111111111111111111; 
assign wn_re[1025] = 26'b11111111111111110000000000; assign wn_im[1025] = 26'b00000000000000000000000011; 
assign wn_re[1026] = 26'b11111111111111110000000000; assign wn_im[1026] = 26'b00000000000000000000000110; 
assign wn_re[1027] = 26'b11111111111111110000000000; assign wn_im[1027] = 26'b00000000000000000000001001; 
assign wn_re[1028] = 26'b11111111111111110000000000; assign wn_im[1028] = 26'b00000000000000000000001100; 
assign wn_re[1029] = 26'b11111111111111110000000000; assign wn_im[1029] = 26'b00000000000000000000001111; 
assign wn_re[1030] = 26'b11111111111111110000000000; assign wn_im[1030] = 26'b00000000000000000000010010; 
assign wn_re[1031] = 26'b11111111111111110000000000; assign wn_im[1031] = 26'b00000000000000000000010101; 
assign wn_re[1032] = 26'b11111111111111110000000000; assign wn_im[1032] = 26'b00000000000000000000011001; 
assign wn_re[1033] = 26'b11111111111111110000000000; assign wn_im[1033] = 26'b00000000000000000000011100; 
assign wn_re[1034] = 26'b11111111111111110000000000; assign wn_im[1034] = 26'b00000000000000000000011111; 
assign wn_re[1035] = 26'b11111111111111110000000000; assign wn_im[1035] = 26'b00000000000000000000100010; 
assign wn_re[1036] = 26'b11111111111111110000000000; assign wn_im[1036] = 26'b00000000000000000000100101; 
assign wn_re[1037] = 26'b11111111111111110000000000; assign wn_im[1037] = 26'b00000000000000000000101000; 
assign wn_re[1038] = 26'b11111111111111110000000000; assign wn_im[1038] = 26'b00000000000000000000101011; 
assign wn_re[1039] = 26'b11111111111111110000000001; assign wn_im[1039] = 26'b00000000000000000000101111; 
assign wn_re[1040] = 26'b11111111111111110000000001; assign wn_im[1040] = 26'b00000000000000000000110010; 
assign wn_re[1041] = 26'b11111111111111110000000001; assign wn_im[1041] = 26'b00000000000000000000110101; 
assign wn_re[1042] = 26'b11111111111111110000000001; assign wn_im[1042] = 26'b00000000000000000000111000; 
assign wn_re[1043] = 26'b11111111111111110000000001; assign wn_im[1043] = 26'b00000000000000000000111011; 
assign wn_re[1044] = 26'b11111111111111110000000001; assign wn_im[1044] = 26'b00000000000000000000111110; 
assign wn_re[1045] = 26'b11111111111111110000000010; assign wn_im[1045] = 26'b00000000000000000001000001; 
assign wn_re[1046] = 26'b11111111111111110000000010; assign wn_im[1046] = 26'b00000000000000000001000101; 
assign wn_re[1047] = 26'b11111111111111110000000010; assign wn_im[1047] = 26'b00000000000000000001001000; 
assign wn_re[1048] = 26'b11111111111111110000000010; assign wn_im[1048] = 26'b00000000000000000001001011; 
assign wn_re[1049] = 26'b11111111111111110000000011; assign wn_im[1049] = 26'b00000000000000000001001110; 
assign wn_re[1050] = 26'b11111111111111110000000011; assign wn_im[1050] = 26'b00000000000000000001010001; 
assign wn_re[1051] = 26'b11111111111111110000000011; assign wn_im[1051] = 26'b00000000000000000001010100; 
assign wn_re[1052] = 26'b11111111111111110000000011; assign wn_im[1052] = 26'b00000000000000000001010111; 
assign wn_re[1053] = 26'b11111111111111110000000100; assign wn_im[1053] = 26'b00000000000000000001011010; 
assign wn_re[1054] = 26'b11111111111111110000000100; assign wn_im[1054] = 26'b00000000000000000001011110; 
assign wn_re[1055] = 26'b11111111111111110000000100; assign wn_im[1055] = 26'b00000000000000000001100001; 
assign wn_re[1056] = 26'b11111111111111110000000100; assign wn_im[1056] = 26'b00000000000000000001100100; 
assign wn_re[1057] = 26'b11111111111111110000000101; assign wn_im[1057] = 26'b00000000000000000001100111; 
assign wn_re[1058] = 26'b11111111111111110000000101; assign wn_im[1058] = 26'b00000000000000000001101010; 
assign wn_re[1059] = 26'b11111111111111110000000101; assign wn_im[1059] = 26'b00000000000000000001101101; 
assign wn_re[1060] = 26'b11111111111111110000000110; assign wn_im[1060] = 26'b00000000000000000001110000; 
assign wn_re[1061] = 26'b11111111111111110000000110; assign wn_im[1061] = 26'b00000000000000000001110011; 
assign wn_re[1062] = 26'b11111111111111110000000110; assign wn_im[1062] = 26'b00000000000000000001110111; 
assign wn_re[1063] = 26'b11111111111111110000000111; assign wn_im[1063] = 26'b00000000000000000001111010; 
assign wn_re[1064] = 26'b11111111111111110000000111; assign wn_im[1064] = 26'b00000000000000000001111101; 
assign wn_re[1065] = 26'b11111111111111110000001000; assign wn_im[1065] = 26'b00000000000000000010000000; 
assign wn_re[1066] = 26'b11111111111111110000001000; assign wn_im[1066] = 26'b00000000000000000010000011; 
assign wn_re[1067] = 26'b11111111111111110000001000; assign wn_im[1067] = 26'b00000000000000000010000110; 
assign wn_re[1068] = 26'b11111111111111110000001001; assign wn_im[1068] = 26'b00000000000000000010001001; 
assign wn_re[1069] = 26'b11111111111111110000001001; assign wn_im[1069] = 26'b00000000000000000010001100; 
assign wn_re[1070] = 26'b11111111111111110000001010; assign wn_im[1070] = 26'b00000000000000000010010000; 
assign wn_re[1071] = 26'b11111111111111110000001010; assign wn_im[1071] = 26'b00000000000000000010010011; 
assign wn_re[1072] = 26'b11111111111111110000001011; assign wn_im[1072] = 26'b00000000000000000010010110; 
assign wn_re[1073] = 26'b11111111111111110000001011; assign wn_im[1073] = 26'b00000000000000000010011001; 
assign wn_re[1074] = 26'b11111111111111110000001100; assign wn_im[1074] = 26'b00000000000000000010011100; 
assign wn_re[1075] = 26'b11111111111111110000001100; assign wn_im[1075] = 26'b00000000000000000010011111; 
assign wn_re[1076] = 26'b11111111111111110000001101; assign wn_im[1076] = 26'b00000000000000000010100010; 
assign wn_re[1077] = 26'b11111111111111110000001101; assign wn_im[1077] = 26'b00000000000000000010100101; 
assign wn_re[1078] = 26'b11111111111111110000001110; assign wn_im[1078] = 26'b00000000000000000010101000; 
assign wn_re[1079] = 26'b11111111111111110000001110; assign wn_im[1079] = 26'b00000000000000000010101011; 
assign wn_re[1080] = 26'b11111111111111110000001111; assign wn_im[1080] = 26'b00000000000000000010101111; 
assign wn_re[1081] = 26'b11111111111111110000001111; assign wn_im[1081] = 26'b00000000000000000010110010; 
assign wn_re[1082] = 26'b11111111111111110000010000; assign wn_im[1082] = 26'b00000000000000000010110101; 
assign wn_re[1083] = 26'b11111111111111110000010000; assign wn_im[1083] = 26'b00000000000000000010111000; 
assign wn_re[1084] = 26'b11111111111111110000010001; assign wn_im[1084] = 26'b00000000000000000010111011; 
assign wn_re[1085] = 26'b11111111111111110000010001; assign wn_im[1085] = 26'b00000000000000000010111110; 
assign wn_re[1086] = 26'b11111111111111110000010010; assign wn_im[1086] = 26'b00000000000000000011000001; 
assign wn_re[1087] = 26'b11111111111111110000010011; assign wn_im[1087] = 26'b00000000000000000011000100; 
assign wn_re[1088] = 26'b11111111111111110000010011; assign wn_im[1088] = 26'b00000000000000000011000111; 
assign wn_re[1089] = 26'b11111111111111110000010100; assign wn_im[1089] = 26'b00000000000000000011001010; 
assign wn_re[1090] = 26'b11111111111111110000010100; assign wn_im[1090] = 26'b00000000000000000011001101; 
assign wn_re[1091] = 26'b11111111111111110000010101; assign wn_im[1091] = 26'b00000000000000000011010001; 
assign wn_re[1092] = 26'b11111111111111110000010110; assign wn_im[1092] = 26'b00000000000000000011010100; 
assign wn_re[1093] = 26'b11111111111111110000010110; assign wn_im[1093] = 26'b00000000000000000011010111; 
assign wn_re[1094] = 26'b11111111111111110000010111; assign wn_im[1094] = 26'b00000000000000000011011010; 
assign wn_re[1095] = 26'b11111111111111110000011000; assign wn_im[1095] = 26'b00000000000000000011011101; 
assign wn_re[1096] = 26'b11111111111111110000011000; assign wn_im[1096] = 26'b00000000000000000011100000; 
assign wn_re[1097] = 26'b11111111111111110000011001; assign wn_im[1097] = 26'b00000000000000000011100011; 
assign wn_re[1098] = 26'b11111111111111110000011010; assign wn_im[1098] = 26'b00000000000000000011100110; 
assign wn_re[1099] = 26'b11111111111111110000011010; assign wn_im[1099] = 26'b00000000000000000011101001; 
assign wn_re[1100] = 26'b11111111111111110000011011; assign wn_im[1100] = 26'b00000000000000000011101100; 
assign wn_re[1101] = 26'b11111111111111110000011100; assign wn_im[1101] = 26'b00000000000000000011101111; 
assign wn_re[1102] = 26'b11111111111111110000011101; assign wn_im[1102] = 26'b00000000000000000011110010; 
assign wn_re[1103] = 26'b11111111111111110000011101; assign wn_im[1103] = 26'b00000000000000000011110101; 
assign wn_re[1104] = 26'b11111111111111110000011110; assign wn_im[1104] = 26'b00000000000000000011111000; 
assign wn_re[1105] = 26'b11111111111111110000011111; assign wn_im[1105] = 26'b00000000000000000011111011; 
assign wn_re[1106] = 26'b11111111111111110000100000; assign wn_im[1106] = 26'b00000000000000000011111110; 
assign wn_re[1107] = 26'b11111111111111110000100001; assign wn_im[1107] = 26'b00000000000000000100000001; 
assign wn_re[1108] = 26'b11111111111111110000100001; assign wn_im[1108] = 26'b00000000000000000100000100; 
assign wn_re[1109] = 26'b11111111111111110000100010; assign wn_im[1109] = 26'b00000000000000000100001000; 
assign wn_re[1110] = 26'b11111111111111110000100011; assign wn_im[1110] = 26'b00000000000000000100001011; 
assign wn_re[1111] = 26'b11111111111111110000100100; assign wn_im[1111] = 26'b00000000000000000100001110; 
assign wn_re[1112] = 26'b11111111111111110000100101; assign wn_im[1112] = 26'b00000000000000000100010001; 
assign wn_re[1113] = 26'b11111111111111110000100101; assign wn_im[1113] = 26'b00000000000000000100010100; 
assign wn_re[1114] = 26'b11111111111111110000100110; assign wn_im[1114] = 26'b00000000000000000100010111; 
assign wn_re[1115] = 26'b11111111111111110000100111; assign wn_im[1115] = 26'b00000000000000000100011010; 
assign wn_re[1116] = 26'b11111111111111110000101000; assign wn_im[1116] = 26'b00000000000000000100011101; 
assign wn_re[1117] = 26'b11111111111111110000101001; assign wn_im[1117] = 26'b00000000000000000100100000; 
assign wn_re[1118] = 26'b11111111111111110000101010; assign wn_im[1118] = 26'b00000000000000000100100011; 
assign wn_re[1119] = 26'b11111111111111110000101011; assign wn_im[1119] = 26'b00000000000000000100100110; 
assign wn_re[1120] = 26'b11111111111111110000101100; assign wn_im[1120] = 26'b00000000000000000100101001; 
assign wn_re[1121] = 26'b11111111111111110000101101; assign wn_im[1121] = 26'b00000000000000000100101100; 
assign wn_re[1122] = 26'b11111111111111110000101101; assign wn_im[1122] = 26'b00000000000000000100101111; 
assign wn_re[1123] = 26'b11111111111111110000101110; assign wn_im[1123] = 26'b00000000000000000100110010; 
assign wn_re[1124] = 26'b11111111111111110000101111; assign wn_im[1124] = 26'b00000000000000000100110101; 
assign wn_re[1125] = 26'b11111111111111110000110000; assign wn_im[1125] = 26'b00000000000000000100111000; 
assign wn_re[1126] = 26'b11111111111111110000110001; assign wn_im[1126] = 26'b00000000000000000100111011; 
assign wn_re[1127] = 26'b11111111111111110000110010; assign wn_im[1127] = 26'b00000000000000000100111110; 
assign wn_re[1128] = 26'b11111111111111110000110011; assign wn_im[1128] = 26'b00000000000000000101000001; 
assign wn_re[1129] = 26'b11111111111111110000110100; assign wn_im[1129] = 26'b00000000000000000101000100; 
assign wn_re[1130] = 26'b11111111111111110000110101; assign wn_im[1130] = 26'b00000000000000000101000111; 
assign wn_re[1131] = 26'b11111111111111110000110110; assign wn_im[1131] = 26'b00000000000000000101001010; 
assign wn_re[1132] = 26'b11111111111111110000110111; assign wn_im[1132] = 26'b00000000000000000101001101; 
assign wn_re[1133] = 26'b11111111111111110000111000; assign wn_im[1133] = 26'b00000000000000000101010000; 
assign wn_re[1134] = 26'b11111111111111110000111001; assign wn_im[1134] = 26'b00000000000000000101010011; 
assign wn_re[1135] = 26'b11111111111111110000111010; assign wn_im[1135] = 26'b00000000000000000101010110; 
assign wn_re[1136] = 26'b11111111111111110000111011; assign wn_im[1136] = 26'b00000000000000000101011000; 
assign wn_re[1137] = 26'b11111111111111110000111100; assign wn_im[1137] = 26'b00000000000000000101011011; 
assign wn_re[1138] = 26'b11111111111111110000111101; assign wn_im[1138] = 26'b00000000000000000101011110; 
assign wn_re[1139] = 26'b11111111111111110000111111; assign wn_im[1139] = 26'b00000000000000000101100001; 
assign wn_re[1140] = 26'b11111111111111110001000000; assign wn_im[1140] = 26'b00000000000000000101100100; 
assign wn_re[1141] = 26'b11111111111111110001000001; assign wn_im[1141] = 26'b00000000000000000101100111; 
assign wn_re[1142] = 26'b11111111111111110001000010; assign wn_im[1142] = 26'b00000000000000000101101010; 
assign wn_re[1143] = 26'b11111111111111110001000011; assign wn_im[1143] = 26'b00000000000000000101101101; 
assign wn_re[1144] = 26'b11111111111111110001000100; assign wn_im[1144] = 26'b00000000000000000101110000; 
assign wn_re[1145] = 26'b11111111111111110001000101; assign wn_im[1145] = 26'b00000000000000000101110011; 
assign wn_re[1146] = 26'b11111111111111110001000110; assign wn_im[1146] = 26'b00000000000000000101110110; 
assign wn_re[1147] = 26'b11111111111111110001001000; assign wn_im[1147] = 26'b00000000000000000101111001; 
assign wn_re[1148] = 26'b11111111111111110001001001; assign wn_im[1148] = 26'b00000000000000000101111100; 
assign wn_re[1149] = 26'b11111111111111110001001010; assign wn_im[1149] = 26'b00000000000000000101111111; 
assign wn_re[1150] = 26'b11111111111111110001001011; assign wn_im[1150] = 26'b00000000000000000110000010; 
assign wn_re[1151] = 26'b11111111111111110001001100; assign wn_im[1151] = 26'b00000000000000000110000100; 
assign wn_re[1152] = 26'b11111111111111110001001101; assign wn_im[1152] = 26'b00000000000000000110000111; 
assign wn_re[1153] = 26'b11111111111111110001001111; assign wn_im[1153] = 26'b00000000000000000110001010; 
assign wn_re[1154] = 26'b11111111111111110001010000; assign wn_im[1154] = 26'b00000000000000000110001101; 
assign wn_re[1155] = 26'b11111111111111110001010001; assign wn_im[1155] = 26'b00000000000000000110010000; 
assign wn_re[1156] = 26'b11111111111111110001010010; assign wn_im[1156] = 26'b00000000000000000110010011; 
assign wn_re[1157] = 26'b11111111111111110001010100; assign wn_im[1157] = 26'b00000000000000000110010110; 
assign wn_re[1158] = 26'b11111111111111110001010101; assign wn_im[1158] = 26'b00000000000000000110011001; 
assign wn_re[1159] = 26'b11111111111111110001010110; assign wn_im[1159] = 26'b00000000000000000110011100; 
assign wn_re[1160] = 26'b11111111111111110001010111; assign wn_im[1160] = 26'b00000000000000000110011110; 
assign wn_re[1161] = 26'b11111111111111110001011001; assign wn_im[1161] = 26'b00000000000000000110100001; 
assign wn_re[1162] = 26'b11111111111111110001011010; assign wn_im[1162] = 26'b00000000000000000110100100; 
assign wn_re[1163] = 26'b11111111111111110001011011; assign wn_im[1163] = 26'b00000000000000000110100111; 
assign wn_re[1164] = 26'b11111111111111110001011101; assign wn_im[1164] = 26'b00000000000000000110101010; 
assign wn_re[1165] = 26'b11111111111111110001011110; assign wn_im[1165] = 26'b00000000000000000110101101; 
assign wn_re[1166] = 26'b11111111111111110001011111; assign wn_im[1166] = 26'b00000000000000000110110000; 
assign wn_re[1167] = 26'b11111111111111110001100000; assign wn_im[1167] = 26'b00000000000000000110110010; 
assign wn_re[1168] = 26'b11111111111111110001100010; assign wn_im[1168] = 26'b00000000000000000110110101; 
assign wn_re[1169] = 26'b11111111111111110001100011; assign wn_im[1169] = 26'b00000000000000000110111000; 
assign wn_re[1170] = 26'b11111111111111110001100101; assign wn_im[1170] = 26'b00000000000000000110111011; 
assign wn_re[1171] = 26'b11111111111111110001100110; assign wn_im[1171] = 26'b00000000000000000110111110; 
assign wn_re[1172] = 26'b11111111111111110001100111; assign wn_im[1172] = 26'b00000000000000000111000001; 
assign wn_re[1173] = 26'b11111111111111110001101001; assign wn_im[1173] = 26'b00000000000000000111000011; 
assign wn_re[1174] = 26'b11111111111111110001101010; assign wn_im[1174] = 26'b00000000000000000111000110; 
assign wn_re[1175] = 26'b11111111111111110001101011; assign wn_im[1175] = 26'b00000000000000000111001001; 
assign wn_re[1176] = 26'b11111111111111110001101101; assign wn_im[1176] = 26'b00000000000000000111001100; 
assign wn_re[1177] = 26'b11111111111111110001101110; assign wn_im[1177] = 26'b00000000000000000111001111; 
assign wn_re[1178] = 26'b11111111111111110001110000; assign wn_im[1178] = 26'b00000000000000000111010010; 
assign wn_re[1179] = 26'b11111111111111110001110001; assign wn_im[1179] = 26'b00000000000000000111010100; 
assign wn_re[1180] = 26'b11111111111111110001110011; assign wn_im[1180] = 26'b00000000000000000111010111; 
assign wn_re[1181] = 26'b11111111111111110001110100; assign wn_im[1181] = 26'b00000000000000000111011010; 
assign wn_re[1182] = 26'b11111111111111110001110101; assign wn_im[1182] = 26'b00000000000000000111011101; 
assign wn_re[1183] = 26'b11111111111111110001110111; assign wn_im[1183] = 26'b00000000000000000111011111; 
assign wn_re[1184] = 26'b11111111111111110001111000; assign wn_im[1184] = 26'b00000000000000000111100010; 
assign wn_re[1185] = 26'b11111111111111110001111010; assign wn_im[1185] = 26'b00000000000000000111100101; 
assign wn_re[1186] = 26'b11111111111111110001111011; assign wn_im[1186] = 26'b00000000000000000111101000; 
assign wn_re[1187] = 26'b11111111111111110001111101; assign wn_im[1187] = 26'b00000000000000000111101011; 
assign wn_re[1188] = 26'b11111111111111110001111110; assign wn_im[1188] = 26'b00000000000000000111101101; 
assign wn_re[1189] = 26'b11111111111111110010000000; assign wn_im[1189] = 26'b00000000000000000111110000; 
assign wn_re[1190] = 26'b11111111111111110010000001; assign wn_im[1190] = 26'b00000000000000000111110011; 
assign wn_re[1191] = 26'b11111111111111110010000011; assign wn_im[1191] = 26'b00000000000000000111110101; 
assign wn_re[1192] = 26'b11111111111111110010000101; assign wn_im[1192] = 26'b00000000000000000111111000; 
assign wn_re[1193] = 26'b11111111111111110010000110; assign wn_im[1193] = 26'b00000000000000000111111011; 
assign wn_re[1194] = 26'b11111111111111110010001000; assign wn_im[1194] = 26'b00000000000000000111111110; 
assign wn_re[1195] = 26'b11111111111111110010001001; assign wn_im[1195] = 26'b00000000000000001000000000; 
assign wn_re[1196] = 26'b11111111111111110010001011; assign wn_im[1196] = 26'b00000000000000001000000011; 
assign wn_re[1197] = 26'b11111111111111110010001100; assign wn_im[1197] = 26'b00000000000000001000000110; 
assign wn_re[1198] = 26'b11111111111111110010001110; assign wn_im[1198] = 26'b00000000000000001000001001; 
assign wn_re[1199] = 26'b11111111111111110010010000; assign wn_im[1199] = 26'b00000000000000001000001011; 
assign wn_re[1200] = 26'b11111111111111110010010001; assign wn_im[1200] = 26'b00000000000000001000001110; 
assign wn_re[1201] = 26'b11111111111111110010010011; assign wn_im[1201] = 26'b00000000000000001000010001; 
assign wn_re[1202] = 26'b11111111111111110010010100; assign wn_im[1202] = 26'b00000000000000001000010011; 
assign wn_re[1203] = 26'b11111111111111110010010110; assign wn_im[1203] = 26'b00000000000000001000010110; 
assign wn_re[1204] = 26'b11111111111111110010011000; assign wn_im[1204] = 26'b00000000000000001000011001; 
assign wn_re[1205] = 26'b11111111111111110010011001; assign wn_im[1205] = 26'b00000000000000001000011011; 
assign wn_re[1206] = 26'b11111111111111110010011011; assign wn_im[1206] = 26'b00000000000000001000011110; 
assign wn_re[1207] = 26'b11111111111111110010011101; assign wn_im[1207] = 26'b00000000000000001000100001; 
assign wn_re[1208] = 26'b11111111111111110010011110; assign wn_im[1208] = 26'b00000000000000001000100011; 
assign wn_re[1209] = 26'b11111111111111110010100000; assign wn_im[1209] = 26'b00000000000000001000100110; 
assign wn_re[1210] = 26'b11111111111111110010100010; assign wn_im[1210] = 26'b00000000000000001000101001; 
assign wn_re[1211] = 26'b11111111111111110010100011; assign wn_im[1211] = 26'b00000000000000001000101011; 
assign wn_re[1212] = 26'b11111111111111110010100101; assign wn_im[1212] = 26'b00000000000000001000101110; 
assign wn_re[1213] = 26'b11111111111111110010100111; assign wn_im[1213] = 26'b00000000000000001000110001; 
assign wn_re[1214] = 26'b11111111111111110010101001; assign wn_im[1214] = 26'b00000000000000001000110011; 
assign wn_re[1215] = 26'b11111111111111110010101010; assign wn_im[1215] = 26'b00000000000000001000110110; 
assign wn_re[1216] = 26'b11111111111111110010101100; assign wn_im[1216] = 26'b00000000000000001000111000; 
assign wn_re[1217] = 26'b11111111111111110010101110; assign wn_im[1217] = 26'b00000000000000001000111011; 
assign wn_re[1218] = 26'b11111111111111110010110000; assign wn_im[1218] = 26'b00000000000000001000111110; 
assign wn_re[1219] = 26'b11111111111111110010110001; assign wn_im[1219] = 26'b00000000000000001001000000; 
assign wn_re[1220] = 26'b11111111111111110010110011; assign wn_im[1220] = 26'b00000000000000001001000011; 
assign wn_re[1221] = 26'b11111111111111110010110101; assign wn_im[1221] = 26'b00000000000000001001000101; 
assign wn_re[1222] = 26'b11111111111111110010110111; assign wn_im[1222] = 26'b00000000000000001001001000; 
assign wn_re[1223] = 26'b11111111111111110010111000; assign wn_im[1223] = 26'b00000000000000001001001011; 
assign wn_re[1224] = 26'b11111111111111110010111010; assign wn_im[1224] = 26'b00000000000000001001001101; 
assign wn_re[1225] = 26'b11111111111111110010111100; assign wn_im[1225] = 26'b00000000000000001001010000; 
assign wn_re[1226] = 26'b11111111111111110010111110; assign wn_im[1226] = 26'b00000000000000001001010010; 
assign wn_re[1227] = 26'b11111111111111110011000000; assign wn_im[1227] = 26'b00000000000000001001010101; 
assign wn_re[1228] = 26'b11111111111111110011000010; assign wn_im[1228] = 26'b00000000000000001001010111; 
assign wn_re[1229] = 26'b11111111111111110011000011; assign wn_im[1229] = 26'b00000000000000001001011010; 
assign wn_re[1230] = 26'b11111111111111110011000101; assign wn_im[1230] = 26'b00000000000000001001011100; 
assign wn_re[1231] = 26'b11111111111111110011000111; assign wn_im[1231] = 26'b00000000000000001001011111; 
assign wn_re[1232] = 26'b11111111111111110011001001; assign wn_im[1232] = 26'b00000000000000001001100001; 
assign wn_re[1233] = 26'b11111111111111110011001011; assign wn_im[1233] = 26'b00000000000000001001100100; 
assign wn_re[1234] = 26'b11111111111111110011001101; assign wn_im[1234] = 26'b00000000000000001001100111; 
assign wn_re[1235] = 26'b11111111111111110011001111; assign wn_im[1235] = 26'b00000000000000001001101001; 
assign wn_re[1236] = 26'b11111111111111110011010001; assign wn_im[1236] = 26'b00000000000000001001101100; 
assign wn_re[1237] = 26'b11111111111111110011010010; assign wn_im[1237] = 26'b00000000000000001001101110; 
assign wn_re[1238] = 26'b11111111111111110011010100; assign wn_im[1238] = 26'b00000000000000001001110001; 
assign wn_re[1239] = 26'b11111111111111110011010110; assign wn_im[1239] = 26'b00000000000000001001110011; 
assign wn_re[1240] = 26'b11111111111111110011011000; assign wn_im[1240] = 26'b00000000000000001001110101; 
assign wn_re[1241] = 26'b11111111111111110011011010; assign wn_im[1241] = 26'b00000000000000001001111000; 
assign wn_re[1242] = 26'b11111111111111110011011100; assign wn_im[1242] = 26'b00000000000000001001111010; 
assign wn_re[1243] = 26'b11111111111111110011011110; assign wn_im[1243] = 26'b00000000000000001001111101; 
assign wn_re[1244] = 26'b11111111111111110011100000; assign wn_im[1244] = 26'b00000000000000001001111111; 
assign wn_re[1245] = 26'b11111111111111110011100010; assign wn_im[1245] = 26'b00000000000000001010000010; 
assign wn_re[1246] = 26'b11111111111111110011100100; assign wn_im[1246] = 26'b00000000000000001010000100; 
assign wn_re[1247] = 26'b11111111111111110011100110; assign wn_im[1247] = 26'b00000000000000001010000111; 
assign wn_re[1248] = 26'b11111111111111110011101000; assign wn_im[1248] = 26'b00000000000000001010001001; 
assign wn_re[1249] = 26'b11111111111111110011101010; assign wn_im[1249] = 26'b00000000000000001010001100; 
assign wn_re[1250] = 26'b11111111111111110011101100; assign wn_im[1250] = 26'b00000000000000001010001110; 
assign wn_re[1251] = 26'b11111111111111110011101110; assign wn_im[1251] = 26'b00000000000000001010010000; 
assign wn_re[1252] = 26'b11111111111111110011110000; assign wn_im[1252] = 26'b00000000000000001010010011; 
assign wn_re[1253] = 26'b11111111111111110011110010; assign wn_im[1253] = 26'b00000000000000001010010101; 
assign wn_re[1254] = 26'b11111111111111110011110100; assign wn_im[1254] = 26'b00000000000000001010011000; 
assign wn_re[1255] = 26'b11111111111111110011110110; assign wn_im[1255] = 26'b00000000000000001010011010; 
assign wn_re[1256] = 26'b11111111111111110011111000; assign wn_im[1256] = 26'b00000000000000001010011100; 
assign wn_re[1257] = 26'b11111111111111110011111010; assign wn_im[1257] = 26'b00000000000000001010011111; 
assign wn_re[1258] = 26'b11111111111111110011111100; assign wn_im[1258] = 26'b00000000000000001010100001; 
assign wn_re[1259] = 26'b11111111111111110011111110; assign wn_im[1259] = 26'b00000000000000001010100011; 
assign wn_re[1260] = 26'b11111111111111110100000000; assign wn_im[1260] = 26'b00000000000000001010100110; 
assign wn_re[1261] = 26'b11111111111111110100000010; assign wn_im[1261] = 26'b00000000000000001010101000; 
assign wn_re[1262] = 26'b11111111111111110100000101; assign wn_im[1262] = 26'b00000000000000001010101011; 
assign wn_re[1263] = 26'b11111111111111110100000111; assign wn_im[1263] = 26'b00000000000000001010101101; 
assign wn_re[1264] = 26'b11111111111111110100001001; assign wn_im[1264] = 26'b00000000000000001010101111; 
assign wn_re[1265] = 26'b11111111111111110100001011; assign wn_im[1265] = 26'b00000000000000001010110010; 
assign wn_re[1266] = 26'b11111111111111110100001101; assign wn_im[1266] = 26'b00000000000000001010110100; 
assign wn_re[1267] = 26'b11111111111111110100001111; assign wn_im[1267] = 26'b00000000000000001010110110; 
assign wn_re[1268] = 26'b11111111111111110100010001; assign wn_im[1268] = 26'b00000000000000001010111000; 
assign wn_re[1269] = 26'b11111111111111110100010011; assign wn_im[1269] = 26'b00000000000000001010111011; 
assign wn_re[1270] = 26'b11111111111111110100010110; assign wn_im[1270] = 26'b00000000000000001010111101; 
assign wn_re[1271] = 26'b11111111111111110100011000; assign wn_im[1271] = 26'b00000000000000001010111111; 
assign wn_re[1272] = 26'b11111111111111110100011010; assign wn_im[1272] = 26'b00000000000000001011000010; 
assign wn_re[1273] = 26'b11111111111111110100011100; assign wn_im[1273] = 26'b00000000000000001011000100; 
assign wn_re[1274] = 26'b11111111111111110100011110; assign wn_im[1274] = 26'b00000000000000001011000110; 
assign wn_re[1275] = 26'b11111111111111110100100000; assign wn_im[1275] = 26'b00000000000000001011001000; 
assign wn_re[1276] = 26'b11111111111111110100100011; assign wn_im[1276] = 26'b00000000000000001011001011; 
assign wn_re[1277] = 26'b11111111111111110100100101; assign wn_im[1277] = 26'b00000000000000001011001101; 
assign wn_re[1278] = 26'b11111111111111110100100111; assign wn_im[1278] = 26'b00000000000000001011001111; 
assign wn_re[1279] = 26'b11111111111111110100101001; assign wn_im[1279] = 26'b00000000000000001011010001; 
assign wn_re[1280] = 26'b11111111111111110100101011; assign wn_im[1280] = 26'b00000000000000001011010100; 
assign wn_re[1281] = 26'b11111111111111110100101110; assign wn_im[1281] = 26'b00000000000000001011010110; 
assign wn_re[1282] = 26'b11111111111111110100110000; assign wn_im[1282] = 26'b00000000000000001011011000; 
assign wn_re[1283] = 26'b11111111111111110100110010; assign wn_im[1283] = 26'b00000000000000001011011010; 
assign wn_re[1284] = 26'b11111111111111110100110100; assign wn_im[1284] = 26'b00000000000000001011011100; 
assign wn_re[1285] = 26'b11111111111111110100110111; assign wn_im[1285] = 26'b00000000000000001011011111; 
assign wn_re[1286] = 26'b11111111111111110100111001; assign wn_im[1286] = 26'b00000000000000001011100001; 
assign wn_re[1287] = 26'b11111111111111110100111011; assign wn_im[1287] = 26'b00000000000000001011100011; 
assign wn_re[1288] = 26'b11111111111111110100111101; assign wn_im[1288] = 26'b00000000000000001011100101; 
assign wn_re[1289] = 26'b11111111111111110101000000; assign wn_im[1289] = 26'b00000000000000001011100111; 
assign wn_re[1290] = 26'b11111111111111110101000010; assign wn_im[1290] = 26'b00000000000000001011101001; 
assign wn_re[1291] = 26'b11111111111111110101000100; assign wn_im[1291] = 26'b00000000000000001011101100; 
assign wn_re[1292] = 26'b11111111111111110101000111; assign wn_im[1292] = 26'b00000000000000001011101110; 
assign wn_re[1293] = 26'b11111111111111110101001001; assign wn_im[1293] = 26'b00000000000000001011110000; 
assign wn_re[1294] = 26'b11111111111111110101001011; assign wn_im[1294] = 26'b00000000000000001011110010; 
assign wn_re[1295] = 26'b11111111111111110101001101; assign wn_im[1295] = 26'b00000000000000001011110100; 
assign wn_re[1296] = 26'b11111111111111110101010000; assign wn_im[1296] = 26'b00000000000000001011110110; 
assign wn_re[1297] = 26'b11111111111111110101010010; assign wn_im[1297] = 26'b00000000000000001011111000; 
assign wn_re[1298] = 26'b11111111111111110101010100; assign wn_im[1298] = 26'b00000000000000001011111010; 
assign wn_re[1299] = 26'b11111111111111110101010111; assign wn_im[1299] = 26'b00000000000000001011111101; 
assign wn_re[1300] = 26'b11111111111111110101011001; assign wn_im[1300] = 26'b00000000000000001011111111; 
assign wn_re[1301] = 26'b11111111111111110101011100; assign wn_im[1301] = 26'b00000000000000001100000001; 
assign wn_re[1302] = 26'b11111111111111110101011110; assign wn_im[1302] = 26'b00000000000000001100000011; 
assign wn_re[1303] = 26'b11111111111111110101100000; assign wn_im[1303] = 26'b00000000000000001100000101; 
assign wn_re[1304] = 26'b11111111111111110101100011; assign wn_im[1304] = 26'b00000000000000001100000111; 
assign wn_re[1305] = 26'b11111111111111110101100101; assign wn_im[1305] = 26'b00000000000000001100001001; 
assign wn_re[1306] = 26'b11111111111111110101100111; assign wn_im[1306] = 26'b00000000000000001100001011; 
assign wn_re[1307] = 26'b11111111111111110101101010; assign wn_im[1307] = 26'b00000000000000001100001101; 
assign wn_re[1308] = 26'b11111111111111110101101100; assign wn_im[1308] = 26'b00000000000000001100001111; 
assign wn_re[1309] = 26'b11111111111111110101101111; assign wn_im[1309] = 26'b00000000000000001100010001; 
assign wn_re[1310] = 26'b11111111111111110101110001; assign wn_im[1310] = 26'b00000000000000001100010011; 
assign wn_re[1311] = 26'b11111111111111110101110011; assign wn_im[1311] = 26'b00000000000000001100010101; 
assign wn_re[1312] = 26'b11111111111111110101110110; assign wn_im[1312] = 26'b00000000000000001100010111; 
assign wn_re[1313] = 26'b11111111111111110101111000; assign wn_im[1313] = 26'b00000000000000001100011001; 
assign wn_re[1314] = 26'b11111111111111110101111011; assign wn_im[1314] = 26'b00000000000000001100011011; 
assign wn_re[1315] = 26'b11111111111111110101111101; assign wn_im[1315] = 26'b00000000000000001100011101; 
assign wn_re[1316] = 26'b11111111111111110110000000; assign wn_im[1316] = 26'b00000000000000001100011111; 
assign wn_re[1317] = 26'b11111111111111110110000010; assign wn_im[1317] = 26'b00000000000000001100100001; 
assign wn_re[1318] = 26'b11111111111111110110000101; assign wn_im[1318] = 26'b00000000000000001100100011; 
assign wn_re[1319] = 26'b11111111111111110110000111; assign wn_im[1319] = 26'b00000000000000001100100101; 
assign wn_re[1320] = 26'b11111111111111110110001010; assign wn_im[1320] = 26'b00000000000000001100100111; 
assign wn_re[1321] = 26'b11111111111111110110001100; assign wn_im[1321] = 26'b00000000000000001100101001; 
assign wn_re[1322] = 26'b11111111111111110110001110; assign wn_im[1322] = 26'b00000000000000001100101011; 
assign wn_re[1323] = 26'b11111111111111110110010001; assign wn_im[1323] = 26'b00000000000000001100101101; 
assign wn_re[1324] = 26'b11111111111111110110010011; assign wn_im[1324] = 26'b00000000000000001100101110; 
assign wn_re[1325] = 26'b11111111111111110110010110; assign wn_im[1325] = 26'b00000000000000001100110000; 
assign wn_re[1326] = 26'b11111111111111110110011000; assign wn_im[1326] = 26'b00000000000000001100110010; 
assign wn_re[1327] = 26'b11111111111111110110011011; assign wn_im[1327] = 26'b00000000000000001100110100; 
assign wn_re[1328] = 26'b11111111111111110110011110; assign wn_im[1328] = 26'b00000000000000001100110110; 
assign wn_re[1329] = 26'b11111111111111110110100000; assign wn_im[1329] = 26'b00000000000000001100111000; 
assign wn_re[1330] = 26'b11111111111111110110100011; assign wn_im[1330] = 26'b00000000000000001100111010; 
assign wn_re[1331] = 26'b11111111111111110110100101; assign wn_im[1331] = 26'b00000000000000001100111100; 
assign wn_re[1332] = 26'b11111111111111110110101000; assign wn_im[1332] = 26'b00000000000000001100111101; 
assign wn_re[1333] = 26'b11111111111111110110101010; assign wn_im[1333] = 26'b00000000000000001100111111; 
assign wn_re[1334] = 26'b11111111111111110110101101; assign wn_im[1334] = 26'b00000000000000001101000001; 
assign wn_re[1335] = 26'b11111111111111110110101111; assign wn_im[1335] = 26'b00000000000000001101000011; 
assign wn_re[1336] = 26'b11111111111111110110110010; assign wn_im[1336] = 26'b00000000000000001101000101; 
assign wn_re[1337] = 26'b11111111111111110110110100; assign wn_im[1337] = 26'b00000000000000001101000111; 
assign wn_re[1338] = 26'b11111111111111110110110111; assign wn_im[1338] = 26'b00000000000000001101001000; 
assign wn_re[1339] = 26'b11111111111111110110111010; assign wn_im[1339] = 26'b00000000000000001101001010; 
assign wn_re[1340] = 26'b11111111111111110110111100; assign wn_im[1340] = 26'b00000000000000001101001100; 
assign wn_re[1341] = 26'b11111111111111110110111111; assign wn_im[1341] = 26'b00000000000000001101001110; 
assign wn_re[1342] = 26'b11111111111111110111000001; assign wn_im[1342] = 26'b00000000000000001101001111; 
assign wn_re[1343] = 26'b11111111111111110111000100; assign wn_im[1343] = 26'b00000000000000001101010001; 
assign wn_re[1344] = 26'b11111111111111110111000111; assign wn_im[1344] = 26'b00000000000000001101010011; 
assign wn_re[1345] = 26'b11111111111111110111001001; assign wn_im[1345] = 26'b00000000000000001101010101; 
assign wn_re[1346] = 26'b11111111111111110111001100; assign wn_im[1346] = 26'b00000000000000001101010110; 
assign wn_re[1347] = 26'b11111111111111110111001110; assign wn_im[1347] = 26'b00000000000000001101011000; 
assign wn_re[1348] = 26'b11111111111111110111010001; assign wn_im[1348] = 26'b00000000000000001101011010; 
assign wn_re[1349] = 26'b11111111111111110111010100; assign wn_im[1349] = 26'b00000000000000001101011100; 
assign wn_re[1350] = 26'b11111111111111110111010110; assign wn_im[1350] = 26'b00000000000000001101011101; 
assign wn_re[1351] = 26'b11111111111111110111011001; assign wn_im[1351] = 26'b00000000000000001101011111; 
assign wn_re[1352] = 26'b11111111111111110111011100; assign wn_im[1352] = 26'b00000000000000001101100001; 
assign wn_re[1353] = 26'b11111111111111110111011110; assign wn_im[1353] = 26'b00000000000000001101100010; 
assign wn_re[1354] = 26'b11111111111111110111100001; assign wn_im[1354] = 26'b00000000000000001101100100; 
assign wn_re[1355] = 26'b11111111111111110111100100; assign wn_im[1355] = 26'b00000000000000001101100110; 
assign wn_re[1356] = 26'b11111111111111110111100110; assign wn_im[1356] = 26'b00000000000000001101100111; 
assign wn_re[1357] = 26'b11111111111111110111101001; assign wn_im[1357] = 26'b00000000000000001101101001; 
assign wn_re[1358] = 26'b11111111111111110111101100; assign wn_im[1358] = 26'b00000000000000001101101011; 
assign wn_re[1359] = 26'b11111111111111110111101110; assign wn_im[1359] = 26'b00000000000000001101101100; 
assign wn_re[1360] = 26'b11111111111111110111110001; assign wn_im[1360] = 26'b00000000000000001101101110; 
assign wn_re[1361] = 26'b11111111111111110111110100; assign wn_im[1361] = 26'b00000000000000001101101111; 
assign wn_re[1362] = 26'b11111111111111110111110110; assign wn_im[1362] = 26'b00000000000000001101110001; 
assign wn_re[1363] = 26'b11111111111111110111111001; assign wn_im[1363] = 26'b00000000000000001101110011; 
assign wn_re[1364] = 26'b11111111111111110111111100; assign wn_im[1364] = 26'b00000000000000001101110100; 
assign wn_re[1365] = 26'b11111111111111110111111111; assign wn_im[1365] = 26'b00000000000000001101110110; 
assign wn_re[1366] = 26'b11111111111111111000000001; assign wn_im[1366] = 26'b00000000000000001101110111; 
assign wn_re[1367] = 26'b11111111111111111000000100; assign wn_im[1367] = 26'b00000000000000001101111001; 
assign wn_re[1368] = 26'b11111111111111111000000111; assign wn_im[1368] = 26'b00000000000000001101111010; 
assign wn_re[1369] = 26'b11111111111111111000001010; assign wn_im[1369] = 26'b00000000000000001101111100; 
assign wn_re[1370] = 26'b11111111111111111000001100; assign wn_im[1370] = 26'b00000000000000001101111110; 
assign wn_re[1371] = 26'b11111111111111111000001111; assign wn_im[1371] = 26'b00000000000000001101111111; 
assign wn_re[1372] = 26'b11111111111111111000010010; assign wn_im[1372] = 26'b00000000000000001110000001; 
assign wn_re[1373] = 26'b11111111111111111000010100; assign wn_im[1373] = 26'b00000000000000001110000010; 
assign wn_re[1374] = 26'b11111111111111111000010111; assign wn_im[1374] = 26'b00000000000000001110000100; 
assign wn_re[1375] = 26'b11111111111111111000011010; assign wn_im[1375] = 26'b00000000000000001110000101; 
assign wn_re[1376] = 26'b11111111111111111000011101; assign wn_im[1376] = 26'b00000000000000001110000111; 
assign wn_re[1377] = 26'b11111111111111111000100000; assign wn_im[1377] = 26'b00000000000000001110001000; 
assign wn_re[1378] = 26'b11111111111111111000100010; assign wn_im[1378] = 26'b00000000000000001110001010; 
assign wn_re[1379] = 26'b11111111111111111000100101; assign wn_im[1379] = 26'b00000000000000001110001011; 
assign wn_re[1380] = 26'b11111111111111111000101000; assign wn_im[1380] = 26'b00000000000000001110001100; 
assign wn_re[1381] = 26'b11111111111111111000101011; assign wn_im[1381] = 26'b00000000000000001110001110; 
assign wn_re[1382] = 26'b11111111111111111000101101; assign wn_im[1382] = 26'b00000000000000001110001111; 
assign wn_re[1383] = 26'b11111111111111111000110000; assign wn_im[1383] = 26'b00000000000000001110010001; 
assign wn_re[1384] = 26'b11111111111111111000110011; assign wn_im[1384] = 26'b00000000000000001110010010; 
assign wn_re[1385] = 26'b11111111111111111000110110; assign wn_im[1385] = 26'b00000000000000001110010100; 
assign wn_re[1386] = 26'b11111111111111111000111001; assign wn_im[1386] = 26'b00000000000000001110010101; 
assign wn_re[1387] = 26'b11111111111111111000111100; assign wn_im[1387] = 26'b00000000000000001110010110; 
assign wn_re[1388] = 26'b11111111111111111000111110; assign wn_im[1388] = 26'b00000000000000001110011000; 
assign wn_re[1389] = 26'b11111111111111111001000001; assign wn_im[1389] = 26'b00000000000000001110011001; 
assign wn_re[1390] = 26'b11111111111111111001000100; assign wn_im[1390] = 26'b00000000000000001110011010; 
assign wn_re[1391] = 26'b11111111111111111001000111; assign wn_im[1391] = 26'b00000000000000001110011100; 
assign wn_re[1392] = 26'b11111111111111111001001010; assign wn_im[1392] = 26'b00000000000000001110011101; 
assign wn_re[1393] = 26'b11111111111111111001001101; assign wn_im[1393] = 26'b00000000000000001110011111; 
assign wn_re[1394] = 26'b11111111111111111001001111; assign wn_im[1394] = 26'b00000000000000001110100000; 
assign wn_re[1395] = 26'b11111111111111111001010010; assign wn_im[1395] = 26'b00000000000000001110100001; 
assign wn_re[1396] = 26'b11111111111111111001010101; assign wn_im[1396] = 26'b00000000000000001110100010; 
assign wn_re[1397] = 26'b11111111111111111001011000; assign wn_im[1397] = 26'b00000000000000001110100100; 
assign wn_re[1398] = 26'b11111111111111111001011011; assign wn_im[1398] = 26'b00000000000000001110100101; 
assign wn_re[1399] = 26'b11111111111111111001011110; assign wn_im[1399] = 26'b00000000000000001110100110; 
assign wn_re[1400] = 26'b11111111111111111001100001; assign wn_im[1400] = 26'b00000000000000001110101000; 
assign wn_re[1401] = 26'b11111111111111111001100011; assign wn_im[1401] = 26'b00000000000000001110101001; 
assign wn_re[1402] = 26'b11111111111111111001100110; assign wn_im[1402] = 26'b00000000000000001110101010; 
assign wn_re[1403] = 26'b11111111111111111001101001; assign wn_im[1403] = 26'b00000000000000001110101011; 
assign wn_re[1404] = 26'b11111111111111111001101100; assign wn_im[1404] = 26'b00000000000000001110101101; 
assign wn_re[1405] = 26'b11111111111111111001101111; assign wn_im[1405] = 26'b00000000000000001110101110; 
assign wn_re[1406] = 26'b11111111111111111001110010; assign wn_im[1406] = 26'b00000000000000001110101111; 
assign wn_re[1407] = 26'b11111111111111111001110101; assign wn_im[1407] = 26'b00000000000000001110110000; 
assign wn_re[1408] = 26'b11111111111111111001111000; assign wn_im[1408] = 26'b00000000000000001110110010; 
assign wn_re[1409] = 26'b11111111111111111001111011; assign wn_im[1409] = 26'b00000000000000001110110011; 
assign wn_re[1410] = 26'b11111111111111111001111101; assign wn_im[1410] = 26'b00000000000000001110110100; 
assign wn_re[1411] = 26'b11111111111111111010000000; assign wn_im[1411] = 26'b00000000000000001110110101; 
assign wn_re[1412] = 26'b11111111111111111010000011; assign wn_im[1412] = 26'b00000000000000001110110110; 
assign wn_re[1413] = 26'b11111111111111111010000110; assign wn_im[1413] = 26'b00000000000000001110110111; 
assign wn_re[1414] = 26'b11111111111111111010001001; assign wn_im[1414] = 26'b00000000000000001110111001; 
assign wn_re[1415] = 26'b11111111111111111010001100; assign wn_im[1415] = 26'b00000000000000001110111010; 
assign wn_re[1416] = 26'b11111111111111111010001111; assign wn_im[1416] = 26'b00000000000000001110111011; 
assign wn_re[1417] = 26'b11111111111111111010010010; assign wn_im[1417] = 26'b00000000000000001110111100; 
assign wn_re[1418] = 26'b11111111111111111010010101; assign wn_im[1418] = 26'b00000000000000001110111101; 
assign wn_re[1419] = 26'b11111111111111111010011000; assign wn_im[1419] = 26'b00000000000000001110111110; 
assign wn_re[1420] = 26'b11111111111111111010011011; assign wn_im[1420] = 26'b00000000000000001110111111; 
assign wn_re[1421] = 26'b11111111111111111010011110; assign wn_im[1421] = 26'b00000000000000001111000000; 
assign wn_re[1422] = 26'b11111111111111111010100001; assign wn_im[1422] = 26'b00000000000000001111000010; 
assign wn_re[1423] = 26'b11111111111111111010100100; assign wn_im[1423] = 26'b00000000000000001111000011; 
assign wn_re[1424] = 26'b11111111111111111010100111; assign wn_im[1424] = 26'b00000000000000001111000100; 
assign wn_re[1425] = 26'b11111111111111111010101001; assign wn_im[1425] = 26'b00000000000000001111000101; 
assign wn_re[1426] = 26'b11111111111111111010101100; assign wn_im[1426] = 26'b00000000000000001111000110; 
assign wn_re[1427] = 26'b11111111111111111010101111; assign wn_im[1427] = 26'b00000000000000001111000111; 
assign wn_re[1428] = 26'b11111111111111111010110010; assign wn_im[1428] = 26'b00000000000000001111001000; 
assign wn_re[1429] = 26'b11111111111111111010110101; assign wn_im[1429] = 26'b00000000000000001111001001; 
assign wn_re[1430] = 26'b11111111111111111010111000; assign wn_im[1430] = 26'b00000000000000001111001010; 
assign wn_re[1431] = 26'b11111111111111111010111011; assign wn_im[1431] = 26'b00000000000000001111001011; 
assign wn_re[1432] = 26'b11111111111111111010111110; assign wn_im[1432] = 26'b00000000000000001111001100; 
assign wn_re[1433] = 26'b11111111111111111011000001; assign wn_im[1433] = 26'b00000000000000001111001101; 
assign wn_re[1434] = 26'b11111111111111111011000100; assign wn_im[1434] = 26'b00000000000000001111001110; 
assign wn_re[1435] = 26'b11111111111111111011000111; assign wn_im[1435] = 26'b00000000000000001111001111; 
assign wn_re[1436] = 26'b11111111111111111011001010; assign wn_im[1436] = 26'b00000000000000001111010000; 
assign wn_re[1437] = 26'b11111111111111111011001101; assign wn_im[1437] = 26'b00000000000000001111010001; 
assign wn_re[1438] = 26'b11111111111111111011010000; assign wn_im[1438] = 26'b00000000000000001111010010; 
assign wn_re[1439] = 26'b11111111111111111011010011; assign wn_im[1439] = 26'b00000000000000001111010010; 
assign wn_re[1440] = 26'b11111111111111111011010110; assign wn_im[1440] = 26'b00000000000000001111010011; 
assign wn_re[1441] = 26'b11111111111111111011011001; assign wn_im[1441] = 26'b00000000000000001111010100; 
assign wn_re[1442] = 26'b11111111111111111011011100; assign wn_im[1442] = 26'b00000000000000001111010101; 
assign wn_re[1443] = 26'b11111111111111111011011111; assign wn_im[1443] = 26'b00000000000000001111010110; 
assign wn_re[1444] = 26'b11111111111111111011100010; assign wn_im[1444] = 26'b00000000000000001111010111; 
assign wn_re[1445] = 26'b11111111111111111011100101; assign wn_im[1445] = 26'b00000000000000001111011000; 
assign wn_re[1446] = 26'b11111111111111111011101000; assign wn_im[1446] = 26'b00000000000000001111011001; 
assign wn_re[1447] = 26'b11111111111111111011101011; assign wn_im[1447] = 26'b00000000000000001111011010; 
assign wn_re[1448] = 26'b11111111111111111011101110; assign wn_im[1448] = 26'b00000000000000001111011010; 
assign wn_re[1449] = 26'b11111111111111111011110001; assign wn_im[1449] = 26'b00000000000000001111011011; 
assign wn_re[1450] = 26'b11111111111111111011110100; assign wn_im[1450] = 26'b00000000000000001111011100; 
assign wn_re[1451] = 26'b11111111111111111011110111; assign wn_im[1451] = 26'b00000000000000001111011101; 
assign wn_re[1452] = 26'b11111111111111111011111011; assign wn_im[1452] = 26'b00000000000000001111011110; 
assign wn_re[1453] = 26'b11111111111111111011111110; assign wn_im[1453] = 26'b00000000000000001111011110; 
assign wn_re[1454] = 26'b11111111111111111100000001; assign wn_im[1454] = 26'b00000000000000001111011111; 
assign wn_re[1455] = 26'b11111111111111111100000100; assign wn_im[1455] = 26'b00000000000000001111100000; 
assign wn_re[1456] = 26'b11111111111111111100000111; assign wn_im[1456] = 26'b00000000000000001111100001; 
assign wn_re[1457] = 26'b11111111111111111100001010; assign wn_im[1457] = 26'b00000000000000001111100010; 
assign wn_re[1458] = 26'b11111111111111111100001101; assign wn_im[1458] = 26'b00000000000000001111100010; 
assign wn_re[1459] = 26'b11111111111111111100010000; assign wn_im[1459] = 26'b00000000000000001111100011; 
assign wn_re[1460] = 26'b11111111111111111100010011; assign wn_im[1460] = 26'b00000000000000001111100100; 
assign wn_re[1461] = 26'b11111111111111111100010110; assign wn_im[1461] = 26'b00000000000000001111100101; 
assign wn_re[1462] = 26'b11111111111111111100011001; assign wn_im[1462] = 26'b00000000000000001111100101; 
assign wn_re[1463] = 26'b11111111111111111100011100; assign wn_im[1463] = 26'b00000000000000001111100110; 
assign wn_re[1464] = 26'b11111111111111111100011111; assign wn_im[1464] = 26'b00000000000000001111100111; 
assign wn_re[1465] = 26'b11111111111111111100100010; assign wn_im[1465] = 26'b00000000000000001111100111; 
assign wn_re[1466] = 26'b11111111111111111100100101; assign wn_im[1466] = 26'b00000000000000001111101000; 
assign wn_re[1467] = 26'b11111111111111111100101000; assign wn_im[1467] = 26'b00000000000000001111101001; 
assign wn_re[1468] = 26'b11111111111111111100101011; assign wn_im[1468] = 26'b00000000000000001111101001; 
assign wn_re[1469] = 26'b11111111111111111100101110; assign wn_im[1469] = 26'b00000000000000001111101010; 
assign wn_re[1470] = 26'b11111111111111111100110010; assign wn_im[1470] = 26'b00000000000000001111101011; 
assign wn_re[1471] = 26'b11111111111111111100110101; assign wn_im[1471] = 26'b00000000000000001111101011; 
assign wn_re[1472] = 26'b11111111111111111100111000; assign wn_im[1472] = 26'b00000000000000001111101100; 
assign wn_re[1473] = 26'b11111111111111111100111011; assign wn_im[1473] = 26'b00000000000000001111101100; 
assign wn_re[1474] = 26'b11111111111111111100111110; assign wn_im[1474] = 26'b00000000000000001111101101; 
assign wn_re[1475] = 26'b11111111111111111101000001; assign wn_im[1475] = 26'b00000000000000001111101110; 
assign wn_re[1476] = 26'b11111111111111111101000100; assign wn_im[1476] = 26'b00000000000000001111101110; 
assign wn_re[1477] = 26'b11111111111111111101000111; assign wn_im[1477] = 26'b00000000000000001111101111; 
assign wn_re[1478] = 26'b11111111111111111101001010; assign wn_im[1478] = 26'b00000000000000001111101111; 
assign wn_re[1479] = 26'b11111111111111111101001101; assign wn_im[1479] = 26'b00000000000000001111110000; 
assign wn_re[1480] = 26'b11111111111111111101010000; assign wn_im[1480] = 26'b00000000000000001111110000; 
assign wn_re[1481] = 26'b11111111111111111101010100; assign wn_im[1481] = 26'b00000000000000001111110001; 
assign wn_re[1482] = 26'b11111111111111111101010111; assign wn_im[1482] = 26'b00000000000000001111110001; 
assign wn_re[1483] = 26'b11111111111111111101011010; assign wn_im[1483] = 26'b00000000000000001111110010; 
assign wn_re[1484] = 26'b11111111111111111101011101; assign wn_im[1484] = 26'b00000000000000001111110010; 
assign wn_re[1485] = 26'b11111111111111111101100000; assign wn_im[1485] = 26'b00000000000000001111110011; 
assign wn_re[1486] = 26'b11111111111111111101100011; assign wn_im[1486] = 26'b00000000000000001111110011; 
assign wn_re[1487] = 26'b11111111111111111101100110; assign wn_im[1487] = 26'b00000000000000001111110100; 
assign wn_re[1488] = 26'b11111111111111111101101001; assign wn_im[1488] = 26'b00000000000000001111110100; 
assign wn_re[1489] = 26'b11111111111111111101101100; assign wn_im[1489] = 26'b00000000000000001111110101; 
assign wn_re[1490] = 26'b11111111111111111101101111; assign wn_im[1490] = 26'b00000000000000001111110101; 
assign wn_re[1491] = 26'b11111111111111111101110011; assign wn_im[1491] = 26'b00000000000000001111110110; 
assign wn_re[1492] = 26'b11111111111111111101110110; assign wn_im[1492] = 26'b00000000000000001111110110; 
assign wn_re[1493] = 26'b11111111111111111101111001; assign wn_im[1493] = 26'b00000000000000001111110111; 
assign wn_re[1494] = 26'b11111111111111111101111100; assign wn_im[1494] = 26'b00000000000000001111110111; 
assign wn_re[1495] = 26'b11111111111111111101111111; assign wn_im[1495] = 26'b00000000000000001111110111; 
assign wn_re[1496] = 26'b11111111111111111110000010; assign wn_im[1496] = 26'b00000000000000001111111000; 
assign wn_re[1497] = 26'b11111111111111111110000101; assign wn_im[1497] = 26'b00000000000000001111111000; 
assign wn_re[1498] = 26'b11111111111111111110001000; assign wn_im[1498] = 26'b00000000000000001111111001; 
assign wn_re[1499] = 26'b11111111111111111110001100; assign wn_im[1499] = 26'b00000000000000001111111001; 
assign wn_re[1500] = 26'b11111111111111111110001111; assign wn_im[1500] = 26'b00000000000000001111111001; 
assign wn_re[1501] = 26'b11111111111111111110010010; assign wn_im[1501] = 26'b00000000000000001111111010; 
assign wn_re[1502] = 26'b11111111111111111110010101; assign wn_im[1502] = 26'b00000000000000001111111010; 
assign wn_re[1503] = 26'b11111111111111111110011000; assign wn_im[1503] = 26'b00000000000000001111111010; 
assign wn_re[1504] = 26'b11111111111111111110011011; assign wn_im[1504] = 26'b00000000000000001111111011; 
assign wn_re[1505] = 26'b11111111111111111110011110; assign wn_im[1505] = 26'b00000000000000001111111011; 
assign wn_re[1506] = 26'b11111111111111111110100001; assign wn_im[1506] = 26'b00000000000000001111111011; 
assign wn_re[1507] = 26'b11111111111111111110100101; assign wn_im[1507] = 26'b00000000000000001111111011; 
assign wn_re[1508] = 26'b11111111111111111110101000; assign wn_im[1508] = 26'b00000000000000001111111100; 
assign wn_re[1509] = 26'b11111111111111111110101011; assign wn_im[1509] = 26'b00000000000000001111111100; 
assign wn_re[1510] = 26'b11111111111111111110101110; assign wn_im[1510] = 26'b00000000000000001111111100; 
assign wn_re[1511] = 26'b11111111111111111110110001; assign wn_im[1511] = 26'b00000000000000001111111100; 
assign wn_re[1512] = 26'b11111111111111111110110100; assign wn_im[1512] = 26'b00000000000000001111111101; 
assign wn_re[1513] = 26'b11111111111111111110110111; assign wn_im[1513] = 26'b00000000000000001111111101; 
assign wn_re[1514] = 26'b11111111111111111110111010; assign wn_im[1514] = 26'b00000000000000001111111101; 
assign wn_re[1515] = 26'b11111111111111111110111110; assign wn_im[1515] = 26'b00000000000000001111111101; 
assign wn_re[1516] = 26'b11111111111111111111000001; assign wn_im[1516] = 26'b00000000000000001111111110; 
assign wn_re[1517] = 26'b11111111111111111111000100; assign wn_im[1517] = 26'b00000000000000001111111110; 
assign wn_re[1518] = 26'b11111111111111111111000111; assign wn_im[1518] = 26'b00000000000000001111111110; 
assign wn_re[1519] = 26'b11111111111111111111001010; assign wn_im[1519] = 26'b00000000000000001111111110; 
assign wn_re[1520] = 26'b11111111111111111111001101; assign wn_im[1520] = 26'b00000000000000001111111110; 
assign wn_re[1521] = 26'b11111111111111111111010000; assign wn_im[1521] = 26'b00000000000000001111111110; 
assign wn_re[1522] = 26'b11111111111111111111010100; assign wn_im[1522] = 26'b00000000000000001111111111; 
assign wn_re[1523] = 26'b11111111111111111111010111; assign wn_im[1523] = 26'b00000000000000001111111111; 
assign wn_re[1524] = 26'b11111111111111111111011010; assign wn_im[1524] = 26'b00000000000000001111111111; 
assign wn_re[1525] = 26'b11111111111111111111011101; assign wn_im[1525] = 26'b00000000000000001111111111; 
assign wn_re[1526] = 26'b11111111111111111111100000; assign wn_im[1526] = 26'b00000000000000001111111111; 
assign wn_re[1527] = 26'b11111111111111111111100011; assign wn_im[1527] = 26'b00000000000000001111111111; 
assign wn_re[1528] = 26'b11111111111111111111100110; assign wn_im[1528] = 26'b00000000000000001111111111; 
assign wn_re[1529] = 26'b11111111111111111111101010; assign wn_im[1529] = 26'b00000000000000001111111111; 
assign wn_re[1530] = 26'b11111111111111111111101101; assign wn_im[1530] = 26'b00000000000000001111111111; 
assign wn_re[1531] = 26'b11111111111111111111110000; assign wn_im[1531] = 26'b00000000000000001111111111; 
assign wn_re[1532] = 26'b11111111111111111111110011; assign wn_im[1532] = 26'b00000000000000001111111111; 
assign wn_re[1533] = 26'b11111111111111111111110110; assign wn_im[1533] = 26'b00000000000000001111111111; 
assign wn_re[1534] = 26'b11111111111111111111111001; assign wn_im[1534] = 26'b00000000000000001111111111; 
assign wn_re[1535] = 26'b11111111111111111111111100; assign wn_im[1535] = 26'b00000000000000001111111111; 
assign wn_re[1536] = 26'b11111111111111111111111111; assign wn_im[1536] = 26'b00000000000000010000000000; 
assign wn_re[1537] = 26'b00000000000000000000000011; assign wn_im[1537] = 26'b00000000000000001111111111; 
assign wn_re[1538] = 26'b00000000000000000000000110; assign wn_im[1538] = 26'b00000000000000001111111111; 
assign wn_re[1539] = 26'b00000000000000000000001001; assign wn_im[1539] = 26'b00000000000000001111111111; 
assign wn_re[1540] = 26'b00000000000000000000001100; assign wn_im[1540] = 26'b00000000000000001111111111; 
assign wn_re[1541] = 26'b00000000000000000000001111; assign wn_im[1541] = 26'b00000000000000001111111111; 
assign wn_re[1542] = 26'b00000000000000000000010010; assign wn_im[1542] = 26'b00000000000000001111111111; 
assign wn_re[1543] = 26'b00000000000000000000010101; assign wn_im[1543] = 26'b00000000000000001111111111; 
assign wn_re[1544] = 26'b00000000000000000000011001; assign wn_im[1544] = 26'b00000000000000001111111111; 
assign wn_re[1545] = 26'b00000000000000000000011100; assign wn_im[1545] = 26'b00000000000000001111111111; 
assign wn_re[1546] = 26'b00000000000000000000011111; assign wn_im[1546] = 26'b00000000000000001111111111; 
assign wn_re[1547] = 26'b00000000000000000000100010; assign wn_im[1547] = 26'b00000000000000001111111111; 
assign wn_re[1548] = 26'b00000000000000000000100101; assign wn_im[1548] = 26'b00000000000000001111111111; 
assign wn_re[1549] = 26'b00000000000000000000101000; assign wn_im[1549] = 26'b00000000000000001111111111; 
assign wn_re[1550] = 26'b00000000000000000000101011; assign wn_im[1550] = 26'b00000000000000001111111111; 
assign wn_re[1551] = 26'b00000000000000000000101111; assign wn_im[1551] = 26'b00000000000000001111111110; 
assign wn_re[1552] = 26'b00000000000000000000110010; assign wn_im[1552] = 26'b00000000000000001111111110; 
assign wn_re[1553] = 26'b00000000000000000000110101; assign wn_im[1553] = 26'b00000000000000001111111110; 
assign wn_re[1554] = 26'b00000000000000000000111000; assign wn_im[1554] = 26'b00000000000000001111111110; 
assign wn_re[1555] = 26'b00000000000000000000111011; assign wn_im[1555] = 26'b00000000000000001111111110; 
assign wn_re[1556] = 26'b00000000000000000000111110; assign wn_im[1556] = 26'b00000000000000001111111110; 
assign wn_re[1557] = 26'b00000000000000000001000001; assign wn_im[1557] = 26'b00000000000000001111111101; 
assign wn_re[1558] = 26'b00000000000000000001000101; assign wn_im[1558] = 26'b00000000000000001111111101; 
assign wn_re[1559] = 26'b00000000000000000001001000; assign wn_im[1559] = 26'b00000000000000001111111101; 
assign wn_re[1560] = 26'b00000000000000000001001011; assign wn_im[1560] = 26'b00000000000000001111111101; 
assign wn_re[1561] = 26'b00000000000000000001001110; assign wn_im[1561] = 26'b00000000000000001111111100; 
assign wn_re[1562] = 26'b00000000000000000001010001; assign wn_im[1562] = 26'b00000000000000001111111100; 
assign wn_re[1563] = 26'b00000000000000000001010100; assign wn_im[1563] = 26'b00000000000000001111111100; 
assign wn_re[1564] = 26'b00000000000000000001010111; assign wn_im[1564] = 26'b00000000000000001111111100; 
assign wn_re[1565] = 26'b00000000000000000001011010; assign wn_im[1565] = 26'b00000000000000001111111011; 
assign wn_re[1566] = 26'b00000000000000000001011110; assign wn_im[1566] = 26'b00000000000000001111111011; 
assign wn_re[1567] = 26'b00000000000000000001100001; assign wn_im[1567] = 26'b00000000000000001111111011; 
assign wn_re[1568] = 26'b00000000000000000001100100; assign wn_im[1568] = 26'b00000000000000001111111011; 
assign wn_re[1569] = 26'b00000000000000000001100111; assign wn_im[1569] = 26'b00000000000000001111111010; 
assign wn_re[1570] = 26'b00000000000000000001101010; assign wn_im[1570] = 26'b00000000000000001111111010; 
assign wn_re[1571] = 26'b00000000000000000001101101; assign wn_im[1571] = 26'b00000000000000001111111010; 
assign wn_re[1572] = 26'b00000000000000000001110000; assign wn_im[1572] = 26'b00000000000000001111111001; 
assign wn_re[1573] = 26'b00000000000000000001110011; assign wn_im[1573] = 26'b00000000000000001111111001; 
assign wn_re[1574] = 26'b00000000000000000001110111; assign wn_im[1574] = 26'b00000000000000001111111001; 
assign wn_re[1575] = 26'b00000000000000000001111010; assign wn_im[1575] = 26'b00000000000000001111111000; 
assign wn_re[1576] = 26'b00000000000000000001111101; assign wn_im[1576] = 26'b00000000000000001111111000; 
assign wn_re[1577] = 26'b00000000000000000010000000; assign wn_im[1577] = 26'b00000000000000001111110111; 
assign wn_re[1578] = 26'b00000000000000000010000011; assign wn_im[1578] = 26'b00000000000000001111110111; 
assign wn_re[1579] = 26'b00000000000000000010000110; assign wn_im[1579] = 26'b00000000000000001111110111; 
assign wn_re[1580] = 26'b00000000000000000010001001; assign wn_im[1580] = 26'b00000000000000001111110110; 
assign wn_re[1581] = 26'b00000000000000000010001100; assign wn_im[1581] = 26'b00000000000000001111110110; 
assign wn_re[1582] = 26'b00000000000000000010010000; assign wn_im[1582] = 26'b00000000000000001111110101; 
assign wn_re[1583] = 26'b00000000000000000010010011; assign wn_im[1583] = 26'b00000000000000001111110101; 
assign wn_re[1584] = 26'b00000000000000000010010110; assign wn_im[1584] = 26'b00000000000000001111110100; 
assign wn_re[1585] = 26'b00000000000000000010011001; assign wn_im[1585] = 26'b00000000000000001111110100; 
assign wn_re[1586] = 26'b00000000000000000010011100; assign wn_im[1586] = 26'b00000000000000001111110011; 
assign wn_re[1587] = 26'b00000000000000000010011111; assign wn_im[1587] = 26'b00000000000000001111110011; 
assign wn_re[1588] = 26'b00000000000000000010100010; assign wn_im[1588] = 26'b00000000000000001111110010; 
assign wn_re[1589] = 26'b00000000000000000010100101; assign wn_im[1589] = 26'b00000000000000001111110010; 
assign wn_re[1590] = 26'b00000000000000000010101000; assign wn_im[1590] = 26'b00000000000000001111110001; 
assign wn_re[1591] = 26'b00000000000000000010101011; assign wn_im[1591] = 26'b00000000000000001111110001; 
assign wn_re[1592] = 26'b00000000000000000010101111; assign wn_im[1592] = 26'b00000000000000001111110000; 
assign wn_re[1593] = 26'b00000000000000000010110010; assign wn_im[1593] = 26'b00000000000000001111110000; 
assign wn_re[1594] = 26'b00000000000000000010110101; assign wn_im[1594] = 26'b00000000000000001111101111; 
assign wn_re[1595] = 26'b00000000000000000010111000; assign wn_im[1595] = 26'b00000000000000001111101111; 
assign wn_re[1596] = 26'b00000000000000000010111011; assign wn_im[1596] = 26'b00000000000000001111101110; 
assign wn_re[1597] = 26'b00000000000000000010111110; assign wn_im[1597] = 26'b00000000000000001111101110; 
assign wn_re[1598] = 26'b00000000000000000011000001; assign wn_im[1598] = 26'b00000000000000001111101101; 
assign wn_re[1599] = 26'b00000000000000000011000100; assign wn_im[1599] = 26'b00000000000000001111101100; 
assign wn_re[1600] = 26'b00000000000000000011000111; assign wn_im[1600] = 26'b00000000000000001111101100; 
assign wn_re[1601] = 26'b00000000000000000011001010; assign wn_im[1601] = 26'b00000000000000001111101011; 
assign wn_re[1602] = 26'b00000000000000000011001101; assign wn_im[1602] = 26'b00000000000000001111101011; 
assign wn_re[1603] = 26'b00000000000000000011010001; assign wn_im[1603] = 26'b00000000000000001111101010; 
assign wn_re[1604] = 26'b00000000000000000011010100; assign wn_im[1604] = 26'b00000000000000001111101001; 
assign wn_re[1605] = 26'b00000000000000000011010111; assign wn_im[1605] = 26'b00000000000000001111101001; 
assign wn_re[1606] = 26'b00000000000000000011011010; assign wn_im[1606] = 26'b00000000000000001111101000; 
assign wn_re[1607] = 26'b00000000000000000011011101; assign wn_im[1607] = 26'b00000000000000001111100111; 
assign wn_re[1608] = 26'b00000000000000000011100000; assign wn_im[1608] = 26'b00000000000000001111100111; 
assign wn_re[1609] = 26'b00000000000000000011100011; assign wn_im[1609] = 26'b00000000000000001111100110; 
assign wn_re[1610] = 26'b00000000000000000011100110; assign wn_im[1610] = 26'b00000000000000001111100101; 
assign wn_re[1611] = 26'b00000000000000000011101001; assign wn_im[1611] = 26'b00000000000000001111100101; 
assign wn_re[1612] = 26'b00000000000000000011101100; assign wn_im[1612] = 26'b00000000000000001111100100; 
assign wn_re[1613] = 26'b00000000000000000011101111; assign wn_im[1613] = 26'b00000000000000001111100011; 
assign wn_re[1614] = 26'b00000000000000000011110010; assign wn_im[1614] = 26'b00000000000000001111100010; 
assign wn_re[1615] = 26'b00000000000000000011110101; assign wn_im[1615] = 26'b00000000000000001111100010; 
assign wn_re[1616] = 26'b00000000000000000011111000; assign wn_im[1616] = 26'b00000000000000001111100001; 
assign wn_re[1617] = 26'b00000000000000000011111011; assign wn_im[1617] = 26'b00000000000000001111100000; 
assign wn_re[1618] = 26'b00000000000000000011111110; assign wn_im[1618] = 26'b00000000000000001111011111; 
assign wn_re[1619] = 26'b00000000000000000100000001; assign wn_im[1619] = 26'b00000000000000001111011110; 
assign wn_re[1620] = 26'b00000000000000000100000100; assign wn_im[1620] = 26'b00000000000000001111011110; 
assign wn_re[1621] = 26'b00000000000000000100001000; assign wn_im[1621] = 26'b00000000000000001111011101; 
assign wn_re[1622] = 26'b00000000000000000100001011; assign wn_im[1622] = 26'b00000000000000001111011100; 
assign wn_re[1623] = 26'b00000000000000000100001110; assign wn_im[1623] = 26'b00000000000000001111011011; 
assign wn_re[1624] = 26'b00000000000000000100010001; assign wn_im[1624] = 26'b00000000000000001111011010; 
assign wn_re[1625] = 26'b00000000000000000100010100; assign wn_im[1625] = 26'b00000000000000001111011010; 
assign wn_re[1626] = 26'b00000000000000000100010111; assign wn_im[1626] = 26'b00000000000000001111011001; 
assign wn_re[1627] = 26'b00000000000000000100011010; assign wn_im[1627] = 26'b00000000000000001111011000; 
assign wn_re[1628] = 26'b00000000000000000100011101; assign wn_im[1628] = 26'b00000000000000001111010111; 
assign wn_re[1629] = 26'b00000000000000000100100000; assign wn_im[1629] = 26'b00000000000000001111010110; 
assign wn_re[1630] = 26'b00000000000000000100100011; assign wn_im[1630] = 26'b00000000000000001111010101; 
assign wn_re[1631] = 26'b00000000000000000100100110; assign wn_im[1631] = 26'b00000000000000001111010100; 
assign wn_re[1632] = 26'b00000000000000000100101001; assign wn_im[1632] = 26'b00000000000000001111010011; 
assign wn_re[1633] = 26'b00000000000000000100101100; assign wn_im[1633] = 26'b00000000000000001111010010; 
assign wn_re[1634] = 26'b00000000000000000100101111; assign wn_im[1634] = 26'b00000000000000001111010010; 
assign wn_re[1635] = 26'b00000000000000000100110010; assign wn_im[1635] = 26'b00000000000000001111010001; 
assign wn_re[1636] = 26'b00000000000000000100110101; assign wn_im[1636] = 26'b00000000000000001111010000; 
assign wn_re[1637] = 26'b00000000000000000100111000; assign wn_im[1637] = 26'b00000000000000001111001111; 
assign wn_re[1638] = 26'b00000000000000000100111011; assign wn_im[1638] = 26'b00000000000000001111001110; 
assign wn_re[1639] = 26'b00000000000000000100111110; assign wn_im[1639] = 26'b00000000000000001111001101; 
assign wn_re[1640] = 26'b00000000000000000101000001; assign wn_im[1640] = 26'b00000000000000001111001100; 
assign wn_re[1641] = 26'b00000000000000000101000100; assign wn_im[1641] = 26'b00000000000000001111001011; 
assign wn_re[1642] = 26'b00000000000000000101000111; assign wn_im[1642] = 26'b00000000000000001111001010; 
assign wn_re[1643] = 26'b00000000000000000101001010; assign wn_im[1643] = 26'b00000000000000001111001001; 
assign wn_re[1644] = 26'b00000000000000000101001101; assign wn_im[1644] = 26'b00000000000000001111001000; 
assign wn_re[1645] = 26'b00000000000000000101010000; assign wn_im[1645] = 26'b00000000000000001111000111; 
assign wn_re[1646] = 26'b00000000000000000101010011; assign wn_im[1646] = 26'b00000000000000001111000110; 
assign wn_re[1647] = 26'b00000000000000000101010110; assign wn_im[1647] = 26'b00000000000000001111000101; 
assign wn_re[1648] = 26'b00000000000000000101011000; assign wn_im[1648] = 26'b00000000000000001111000100; 
assign wn_re[1649] = 26'b00000000000000000101011011; assign wn_im[1649] = 26'b00000000000000001111000011; 
assign wn_re[1650] = 26'b00000000000000000101011110; assign wn_im[1650] = 26'b00000000000000001111000010; 
assign wn_re[1651] = 26'b00000000000000000101100001; assign wn_im[1651] = 26'b00000000000000001111000000; 
assign wn_re[1652] = 26'b00000000000000000101100100; assign wn_im[1652] = 26'b00000000000000001110111111; 
assign wn_re[1653] = 26'b00000000000000000101100111; assign wn_im[1653] = 26'b00000000000000001110111110; 
assign wn_re[1654] = 26'b00000000000000000101101010; assign wn_im[1654] = 26'b00000000000000001110111101; 
assign wn_re[1655] = 26'b00000000000000000101101101; assign wn_im[1655] = 26'b00000000000000001110111100; 
assign wn_re[1656] = 26'b00000000000000000101110000; assign wn_im[1656] = 26'b00000000000000001110111011; 
assign wn_re[1657] = 26'b00000000000000000101110011; assign wn_im[1657] = 26'b00000000000000001110111010; 
assign wn_re[1658] = 26'b00000000000000000101110110; assign wn_im[1658] = 26'b00000000000000001110111001; 
assign wn_re[1659] = 26'b00000000000000000101111001; assign wn_im[1659] = 26'b00000000000000001110110111; 
assign wn_re[1660] = 26'b00000000000000000101111100; assign wn_im[1660] = 26'b00000000000000001110110110; 
assign wn_re[1661] = 26'b00000000000000000101111111; assign wn_im[1661] = 26'b00000000000000001110110101; 
assign wn_re[1662] = 26'b00000000000000000110000010; assign wn_im[1662] = 26'b00000000000000001110110100; 
assign wn_re[1663] = 26'b00000000000000000110000100; assign wn_im[1663] = 26'b00000000000000001110110011; 
assign wn_re[1664] = 26'b00000000000000000110000111; assign wn_im[1664] = 26'b00000000000000001110110010; 
assign wn_re[1665] = 26'b00000000000000000110001010; assign wn_im[1665] = 26'b00000000000000001110110000; 
assign wn_re[1666] = 26'b00000000000000000110001101; assign wn_im[1666] = 26'b00000000000000001110101111; 
assign wn_re[1667] = 26'b00000000000000000110010000; assign wn_im[1667] = 26'b00000000000000001110101110; 
assign wn_re[1668] = 26'b00000000000000000110010011; assign wn_im[1668] = 26'b00000000000000001110101101; 
assign wn_re[1669] = 26'b00000000000000000110010110; assign wn_im[1669] = 26'b00000000000000001110101011; 
assign wn_re[1670] = 26'b00000000000000000110011001; assign wn_im[1670] = 26'b00000000000000001110101010; 
assign wn_re[1671] = 26'b00000000000000000110011100; assign wn_im[1671] = 26'b00000000000000001110101001; 
assign wn_re[1672] = 26'b00000000000000000110011110; assign wn_im[1672] = 26'b00000000000000001110101000; 
assign wn_re[1673] = 26'b00000000000000000110100001; assign wn_im[1673] = 26'b00000000000000001110100110; 
assign wn_re[1674] = 26'b00000000000000000110100100; assign wn_im[1674] = 26'b00000000000000001110100101; 
assign wn_re[1675] = 26'b00000000000000000110100111; assign wn_im[1675] = 26'b00000000000000001110100100; 
assign wn_re[1676] = 26'b00000000000000000110101010; assign wn_im[1676] = 26'b00000000000000001110100010; 
assign wn_re[1677] = 26'b00000000000000000110101101; assign wn_im[1677] = 26'b00000000000000001110100001; 
assign wn_re[1678] = 26'b00000000000000000110110000; assign wn_im[1678] = 26'b00000000000000001110100000; 
assign wn_re[1679] = 26'b00000000000000000110110010; assign wn_im[1679] = 26'b00000000000000001110011111; 
assign wn_re[1680] = 26'b00000000000000000110110101; assign wn_im[1680] = 26'b00000000000000001110011101; 
assign wn_re[1681] = 26'b00000000000000000110111000; assign wn_im[1681] = 26'b00000000000000001110011100; 
assign wn_re[1682] = 26'b00000000000000000110111011; assign wn_im[1682] = 26'b00000000000000001110011010; 
assign wn_re[1683] = 26'b00000000000000000110111110; assign wn_im[1683] = 26'b00000000000000001110011001; 
assign wn_re[1684] = 26'b00000000000000000111000001; assign wn_im[1684] = 26'b00000000000000001110011000; 
assign wn_re[1685] = 26'b00000000000000000111000011; assign wn_im[1685] = 26'b00000000000000001110010110; 
assign wn_re[1686] = 26'b00000000000000000111000110; assign wn_im[1686] = 26'b00000000000000001110010101; 
assign wn_re[1687] = 26'b00000000000000000111001001; assign wn_im[1687] = 26'b00000000000000001110010100; 
assign wn_re[1688] = 26'b00000000000000000111001100; assign wn_im[1688] = 26'b00000000000000001110010010; 
assign wn_re[1689] = 26'b00000000000000000111001111; assign wn_im[1689] = 26'b00000000000000001110010001; 
assign wn_re[1690] = 26'b00000000000000000111010010; assign wn_im[1690] = 26'b00000000000000001110001111; 
assign wn_re[1691] = 26'b00000000000000000111010100; assign wn_im[1691] = 26'b00000000000000001110001110; 
assign wn_re[1692] = 26'b00000000000000000111010111; assign wn_im[1692] = 26'b00000000000000001110001100; 
assign wn_re[1693] = 26'b00000000000000000111011010; assign wn_im[1693] = 26'b00000000000000001110001011; 
assign wn_re[1694] = 26'b00000000000000000111011101; assign wn_im[1694] = 26'b00000000000000001110001010; 
assign wn_re[1695] = 26'b00000000000000000111011111; assign wn_im[1695] = 26'b00000000000000001110001000; 
assign wn_re[1696] = 26'b00000000000000000111100010; assign wn_im[1696] = 26'b00000000000000001110000111; 
assign wn_re[1697] = 26'b00000000000000000111100101; assign wn_im[1697] = 26'b00000000000000001110000101; 
assign wn_re[1698] = 26'b00000000000000000111101000; assign wn_im[1698] = 26'b00000000000000001110000100; 
assign wn_re[1699] = 26'b00000000000000000111101011; assign wn_im[1699] = 26'b00000000000000001110000010; 
assign wn_re[1700] = 26'b00000000000000000111101101; assign wn_im[1700] = 26'b00000000000000001110000001; 
assign wn_re[1701] = 26'b00000000000000000111110000; assign wn_im[1701] = 26'b00000000000000001101111111; 
assign wn_re[1702] = 26'b00000000000000000111110011; assign wn_im[1702] = 26'b00000000000000001101111110; 
assign wn_re[1703] = 26'b00000000000000000111110101; assign wn_im[1703] = 26'b00000000000000001101111100; 
assign wn_re[1704] = 26'b00000000000000000111111000; assign wn_im[1704] = 26'b00000000000000001101111010; 
assign wn_re[1705] = 26'b00000000000000000111111011; assign wn_im[1705] = 26'b00000000000000001101111001; 
assign wn_re[1706] = 26'b00000000000000000111111110; assign wn_im[1706] = 26'b00000000000000001101110111; 
assign wn_re[1707] = 26'b00000000000000001000000000; assign wn_im[1707] = 26'b00000000000000001101110110; 
assign wn_re[1708] = 26'b00000000000000001000000011; assign wn_im[1708] = 26'b00000000000000001101110100; 
assign wn_re[1709] = 26'b00000000000000001000000110; assign wn_im[1709] = 26'b00000000000000001101110011; 
assign wn_re[1710] = 26'b00000000000000001000001001; assign wn_im[1710] = 26'b00000000000000001101110001; 
assign wn_re[1711] = 26'b00000000000000001000001011; assign wn_im[1711] = 26'b00000000000000001101101111; 
assign wn_re[1712] = 26'b00000000000000001000001110; assign wn_im[1712] = 26'b00000000000000001101101110; 
assign wn_re[1713] = 26'b00000000000000001000010001; assign wn_im[1713] = 26'b00000000000000001101101100; 
assign wn_re[1714] = 26'b00000000000000001000010011; assign wn_im[1714] = 26'b00000000000000001101101011; 
assign wn_re[1715] = 26'b00000000000000001000010110; assign wn_im[1715] = 26'b00000000000000001101101001; 
assign wn_re[1716] = 26'b00000000000000001000011001; assign wn_im[1716] = 26'b00000000000000001101100111; 
assign wn_re[1717] = 26'b00000000000000001000011011; assign wn_im[1717] = 26'b00000000000000001101100110; 
assign wn_re[1718] = 26'b00000000000000001000011110; assign wn_im[1718] = 26'b00000000000000001101100100; 
assign wn_re[1719] = 26'b00000000000000001000100001; assign wn_im[1719] = 26'b00000000000000001101100010; 
assign wn_re[1720] = 26'b00000000000000001000100011; assign wn_im[1720] = 26'b00000000000000001101100001; 
assign wn_re[1721] = 26'b00000000000000001000100110; assign wn_im[1721] = 26'b00000000000000001101011111; 
assign wn_re[1722] = 26'b00000000000000001000101001; assign wn_im[1722] = 26'b00000000000000001101011101; 
assign wn_re[1723] = 26'b00000000000000001000101011; assign wn_im[1723] = 26'b00000000000000001101011100; 
assign wn_re[1724] = 26'b00000000000000001000101110; assign wn_im[1724] = 26'b00000000000000001101011010; 
assign wn_re[1725] = 26'b00000000000000001000110001; assign wn_im[1725] = 26'b00000000000000001101011000; 
assign wn_re[1726] = 26'b00000000000000001000110011; assign wn_im[1726] = 26'b00000000000000001101010110; 
assign wn_re[1727] = 26'b00000000000000001000110110; assign wn_im[1727] = 26'b00000000000000001101010101; 
assign wn_re[1728] = 26'b00000000000000001000111000; assign wn_im[1728] = 26'b00000000000000001101010011; 
assign wn_re[1729] = 26'b00000000000000001000111011; assign wn_im[1729] = 26'b00000000000000001101010001; 
assign wn_re[1730] = 26'b00000000000000001000111110; assign wn_im[1730] = 26'b00000000000000001101001111; 
assign wn_re[1731] = 26'b00000000000000001001000000; assign wn_im[1731] = 26'b00000000000000001101001110; 
assign wn_re[1732] = 26'b00000000000000001001000011; assign wn_im[1732] = 26'b00000000000000001101001100; 
assign wn_re[1733] = 26'b00000000000000001001000101; assign wn_im[1733] = 26'b00000000000000001101001010; 
assign wn_re[1734] = 26'b00000000000000001001001000; assign wn_im[1734] = 26'b00000000000000001101001000; 
assign wn_re[1735] = 26'b00000000000000001001001011; assign wn_im[1735] = 26'b00000000000000001101000111; 
assign wn_re[1736] = 26'b00000000000000001001001101; assign wn_im[1736] = 26'b00000000000000001101000101; 
assign wn_re[1737] = 26'b00000000000000001001010000; assign wn_im[1737] = 26'b00000000000000001101000011; 
assign wn_re[1738] = 26'b00000000000000001001010010; assign wn_im[1738] = 26'b00000000000000001101000001; 
assign wn_re[1739] = 26'b00000000000000001001010101; assign wn_im[1739] = 26'b00000000000000001100111111; 
assign wn_re[1740] = 26'b00000000000000001001010111; assign wn_im[1740] = 26'b00000000000000001100111101; 
assign wn_re[1741] = 26'b00000000000000001001011010; assign wn_im[1741] = 26'b00000000000000001100111100; 
assign wn_re[1742] = 26'b00000000000000001001011100; assign wn_im[1742] = 26'b00000000000000001100111010; 
assign wn_re[1743] = 26'b00000000000000001001011111; assign wn_im[1743] = 26'b00000000000000001100111000; 
assign wn_re[1744] = 26'b00000000000000001001100001; assign wn_im[1744] = 26'b00000000000000001100110110; 
assign wn_re[1745] = 26'b00000000000000001001100100; assign wn_im[1745] = 26'b00000000000000001100110100; 
assign wn_re[1746] = 26'b00000000000000001001100111; assign wn_im[1746] = 26'b00000000000000001100110010; 
assign wn_re[1747] = 26'b00000000000000001001101001; assign wn_im[1747] = 26'b00000000000000001100110000; 
assign wn_re[1748] = 26'b00000000000000001001101100; assign wn_im[1748] = 26'b00000000000000001100101110; 
assign wn_re[1749] = 26'b00000000000000001001101110; assign wn_im[1749] = 26'b00000000000000001100101101; 
assign wn_re[1750] = 26'b00000000000000001001110001; assign wn_im[1750] = 26'b00000000000000001100101011; 
assign wn_re[1751] = 26'b00000000000000001001110011; assign wn_im[1751] = 26'b00000000000000001100101001; 
assign wn_re[1752] = 26'b00000000000000001001110101; assign wn_im[1752] = 26'b00000000000000001100100111; 
assign wn_re[1753] = 26'b00000000000000001001111000; assign wn_im[1753] = 26'b00000000000000001100100101; 
assign wn_re[1754] = 26'b00000000000000001001111010; assign wn_im[1754] = 26'b00000000000000001100100011; 
assign wn_re[1755] = 26'b00000000000000001001111101; assign wn_im[1755] = 26'b00000000000000001100100001; 
assign wn_re[1756] = 26'b00000000000000001001111111; assign wn_im[1756] = 26'b00000000000000001100011111; 
assign wn_re[1757] = 26'b00000000000000001010000010; assign wn_im[1757] = 26'b00000000000000001100011101; 
assign wn_re[1758] = 26'b00000000000000001010000100; assign wn_im[1758] = 26'b00000000000000001100011011; 
assign wn_re[1759] = 26'b00000000000000001010000111; assign wn_im[1759] = 26'b00000000000000001100011001; 
assign wn_re[1760] = 26'b00000000000000001010001001; assign wn_im[1760] = 26'b00000000000000001100010111; 
assign wn_re[1761] = 26'b00000000000000001010001100; assign wn_im[1761] = 26'b00000000000000001100010101; 
assign wn_re[1762] = 26'b00000000000000001010001110; assign wn_im[1762] = 26'b00000000000000001100010011; 
assign wn_re[1763] = 26'b00000000000000001010010000; assign wn_im[1763] = 26'b00000000000000001100010001; 
assign wn_re[1764] = 26'b00000000000000001010010011; assign wn_im[1764] = 26'b00000000000000001100001111; 
assign wn_re[1765] = 26'b00000000000000001010010101; assign wn_im[1765] = 26'b00000000000000001100001101; 
assign wn_re[1766] = 26'b00000000000000001010011000; assign wn_im[1766] = 26'b00000000000000001100001011; 
assign wn_re[1767] = 26'b00000000000000001010011010; assign wn_im[1767] = 26'b00000000000000001100001001; 
assign wn_re[1768] = 26'b00000000000000001010011100; assign wn_im[1768] = 26'b00000000000000001100000111; 
assign wn_re[1769] = 26'b00000000000000001010011111; assign wn_im[1769] = 26'b00000000000000001100000101; 
assign wn_re[1770] = 26'b00000000000000001010100001; assign wn_im[1770] = 26'b00000000000000001100000011; 
assign wn_re[1771] = 26'b00000000000000001010100011; assign wn_im[1771] = 26'b00000000000000001100000001; 
assign wn_re[1772] = 26'b00000000000000001010100110; assign wn_im[1772] = 26'b00000000000000001011111111; 
assign wn_re[1773] = 26'b00000000000000001010101000; assign wn_im[1773] = 26'b00000000000000001011111101; 
assign wn_re[1774] = 26'b00000000000000001010101011; assign wn_im[1774] = 26'b00000000000000001011111010; 
assign wn_re[1775] = 26'b00000000000000001010101101; assign wn_im[1775] = 26'b00000000000000001011111000; 
assign wn_re[1776] = 26'b00000000000000001010101111; assign wn_im[1776] = 26'b00000000000000001011110110; 
assign wn_re[1777] = 26'b00000000000000001010110010; assign wn_im[1777] = 26'b00000000000000001011110100; 
assign wn_re[1778] = 26'b00000000000000001010110100; assign wn_im[1778] = 26'b00000000000000001011110010; 
assign wn_re[1779] = 26'b00000000000000001010110110; assign wn_im[1779] = 26'b00000000000000001011110000; 
assign wn_re[1780] = 26'b00000000000000001010111000; assign wn_im[1780] = 26'b00000000000000001011101110; 
assign wn_re[1781] = 26'b00000000000000001010111011; assign wn_im[1781] = 26'b00000000000000001011101100; 
assign wn_re[1782] = 26'b00000000000000001010111101; assign wn_im[1782] = 26'b00000000000000001011101001; 
assign wn_re[1783] = 26'b00000000000000001010111111; assign wn_im[1783] = 26'b00000000000000001011100111; 
assign wn_re[1784] = 26'b00000000000000001011000010; assign wn_im[1784] = 26'b00000000000000001011100101; 
assign wn_re[1785] = 26'b00000000000000001011000100; assign wn_im[1785] = 26'b00000000000000001011100011; 
assign wn_re[1786] = 26'b00000000000000001011000110; assign wn_im[1786] = 26'b00000000000000001011100001; 
assign wn_re[1787] = 26'b00000000000000001011001000; assign wn_im[1787] = 26'b00000000000000001011011111; 
assign wn_re[1788] = 26'b00000000000000001011001011; assign wn_im[1788] = 26'b00000000000000001011011100; 
assign wn_re[1789] = 26'b00000000000000001011001101; assign wn_im[1789] = 26'b00000000000000001011011010; 
assign wn_re[1790] = 26'b00000000000000001011001111; assign wn_im[1790] = 26'b00000000000000001011011000; 
assign wn_re[1791] = 26'b00000000000000001011010001; assign wn_im[1791] = 26'b00000000000000001011010110; 
assign wn_re[1792] = 26'b00000000000000001011010100; assign wn_im[1792] = 26'b00000000000000001011010100; 
assign wn_re[1793] = 26'b00000000000000001011010110; assign wn_im[1793] = 26'b00000000000000001011010001; 
assign wn_re[1794] = 26'b00000000000000001011011000; assign wn_im[1794] = 26'b00000000000000001011001111; 
assign wn_re[1795] = 26'b00000000000000001011011010; assign wn_im[1795] = 26'b00000000000000001011001101; 
assign wn_re[1796] = 26'b00000000000000001011011100; assign wn_im[1796] = 26'b00000000000000001011001011; 
assign wn_re[1797] = 26'b00000000000000001011011111; assign wn_im[1797] = 26'b00000000000000001011001000; 
assign wn_re[1798] = 26'b00000000000000001011100001; assign wn_im[1798] = 26'b00000000000000001011000110; 
assign wn_re[1799] = 26'b00000000000000001011100011; assign wn_im[1799] = 26'b00000000000000001011000100; 
assign wn_re[1800] = 26'b00000000000000001011100101; assign wn_im[1800] = 26'b00000000000000001011000010; 
assign wn_re[1801] = 26'b00000000000000001011100111; assign wn_im[1801] = 26'b00000000000000001010111111; 
assign wn_re[1802] = 26'b00000000000000001011101001; assign wn_im[1802] = 26'b00000000000000001010111101; 
assign wn_re[1803] = 26'b00000000000000001011101100; assign wn_im[1803] = 26'b00000000000000001010111011; 
assign wn_re[1804] = 26'b00000000000000001011101110; assign wn_im[1804] = 26'b00000000000000001010111000; 
assign wn_re[1805] = 26'b00000000000000001011110000; assign wn_im[1805] = 26'b00000000000000001010110110; 
assign wn_re[1806] = 26'b00000000000000001011110010; assign wn_im[1806] = 26'b00000000000000001010110100; 
assign wn_re[1807] = 26'b00000000000000001011110100; assign wn_im[1807] = 26'b00000000000000001010110010; 
assign wn_re[1808] = 26'b00000000000000001011110110; assign wn_im[1808] = 26'b00000000000000001010101111; 
assign wn_re[1809] = 26'b00000000000000001011111000; assign wn_im[1809] = 26'b00000000000000001010101101; 
assign wn_re[1810] = 26'b00000000000000001011111010; assign wn_im[1810] = 26'b00000000000000001010101011; 
assign wn_re[1811] = 26'b00000000000000001011111101; assign wn_im[1811] = 26'b00000000000000001010101000; 
assign wn_re[1812] = 26'b00000000000000001011111111; assign wn_im[1812] = 26'b00000000000000001010100110; 
assign wn_re[1813] = 26'b00000000000000001100000001; assign wn_im[1813] = 26'b00000000000000001010100011; 
assign wn_re[1814] = 26'b00000000000000001100000011; assign wn_im[1814] = 26'b00000000000000001010100001; 
assign wn_re[1815] = 26'b00000000000000001100000101; assign wn_im[1815] = 26'b00000000000000001010011111; 
assign wn_re[1816] = 26'b00000000000000001100000111; assign wn_im[1816] = 26'b00000000000000001010011100; 
assign wn_re[1817] = 26'b00000000000000001100001001; assign wn_im[1817] = 26'b00000000000000001010011010; 
assign wn_re[1818] = 26'b00000000000000001100001011; assign wn_im[1818] = 26'b00000000000000001010011000; 
assign wn_re[1819] = 26'b00000000000000001100001101; assign wn_im[1819] = 26'b00000000000000001010010101; 
assign wn_re[1820] = 26'b00000000000000001100001111; assign wn_im[1820] = 26'b00000000000000001010010011; 
assign wn_re[1821] = 26'b00000000000000001100010001; assign wn_im[1821] = 26'b00000000000000001010010000; 
assign wn_re[1822] = 26'b00000000000000001100010011; assign wn_im[1822] = 26'b00000000000000001010001110; 
assign wn_re[1823] = 26'b00000000000000001100010101; assign wn_im[1823] = 26'b00000000000000001010001100; 
assign wn_re[1824] = 26'b00000000000000001100010111; assign wn_im[1824] = 26'b00000000000000001010001001; 
assign wn_re[1825] = 26'b00000000000000001100011001; assign wn_im[1825] = 26'b00000000000000001010000111; 
assign wn_re[1826] = 26'b00000000000000001100011011; assign wn_im[1826] = 26'b00000000000000001010000100; 
assign wn_re[1827] = 26'b00000000000000001100011101; assign wn_im[1827] = 26'b00000000000000001010000010; 
assign wn_re[1828] = 26'b00000000000000001100011111; assign wn_im[1828] = 26'b00000000000000001001111111; 
assign wn_re[1829] = 26'b00000000000000001100100001; assign wn_im[1829] = 26'b00000000000000001001111101; 
assign wn_re[1830] = 26'b00000000000000001100100011; assign wn_im[1830] = 26'b00000000000000001001111010; 
assign wn_re[1831] = 26'b00000000000000001100100101; assign wn_im[1831] = 26'b00000000000000001001111000; 
assign wn_re[1832] = 26'b00000000000000001100100111; assign wn_im[1832] = 26'b00000000000000001001110101; 
assign wn_re[1833] = 26'b00000000000000001100101001; assign wn_im[1833] = 26'b00000000000000001001110011; 
assign wn_re[1834] = 26'b00000000000000001100101011; assign wn_im[1834] = 26'b00000000000000001001110001; 
assign wn_re[1835] = 26'b00000000000000001100101101; assign wn_im[1835] = 26'b00000000000000001001101110; 
assign wn_re[1836] = 26'b00000000000000001100101110; assign wn_im[1836] = 26'b00000000000000001001101100; 
assign wn_re[1837] = 26'b00000000000000001100110000; assign wn_im[1837] = 26'b00000000000000001001101001; 
assign wn_re[1838] = 26'b00000000000000001100110010; assign wn_im[1838] = 26'b00000000000000001001100111; 
assign wn_re[1839] = 26'b00000000000000001100110100; assign wn_im[1839] = 26'b00000000000000001001100100; 
assign wn_re[1840] = 26'b00000000000000001100110110; assign wn_im[1840] = 26'b00000000000000001001100001; 
assign wn_re[1841] = 26'b00000000000000001100111000; assign wn_im[1841] = 26'b00000000000000001001011111; 
assign wn_re[1842] = 26'b00000000000000001100111010; assign wn_im[1842] = 26'b00000000000000001001011100; 
assign wn_re[1843] = 26'b00000000000000001100111100; assign wn_im[1843] = 26'b00000000000000001001011010; 
assign wn_re[1844] = 26'b00000000000000001100111101; assign wn_im[1844] = 26'b00000000000000001001010111; 
assign wn_re[1845] = 26'b00000000000000001100111111; assign wn_im[1845] = 26'b00000000000000001001010101; 
assign wn_re[1846] = 26'b00000000000000001101000001; assign wn_im[1846] = 26'b00000000000000001001010010; 
assign wn_re[1847] = 26'b00000000000000001101000011; assign wn_im[1847] = 26'b00000000000000001001010000; 
assign wn_re[1848] = 26'b00000000000000001101000101; assign wn_im[1848] = 26'b00000000000000001001001101; 
assign wn_re[1849] = 26'b00000000000000001101000111; assign wn_im[1849] = 26'b00000000000000001001001011; 
assign wn_re[1850] = 26'b00000000000000001101001000; assign wn_im[1850] = 26'b00000000000000001001001000; 
assign wn_re[1851] = 26'b00000000000000001101001010; assign wn_im[1851] = 26'b00000000000000001001000101; 
assign wn_re[1852] = 26'b00000000000000001101001100; assign wn_im[1852] = 26'b00000000000000001001000011; 
assign wn_re[1853] = 26'b00000000000000001101001110; assign wn_im[1853] = 26'b00000000000000001001000000; 
assign wn_re[1854] = 26'b00000000000000001101001111; assign wn_im[1854] = 26'b00000000000000001000111110; 
assign wn_re[1855] = 26'b00000000000000001101010001; assign wn_im[1855] = 26'b00000000000000001000111011; 
assign wn_re[1856] = 26'b00000000000000001101010011; assign wn_im[1856] = 26'b00000000000000001000111000; 
assign wn_re[1857] = 26'b00000000000000001101010101; assign wn_im[1857] = 26'b00000000000000001000110110; 
assign wn_re[1858] = 26'b00000000000000001101010110; assign wn_im[1858] = 26'b00000000000000001000110011; 
assign wn_re[1859] = 26'b00000000000000001101011000; assign wn_im[1859] = 26'b00000000000000001000110001; 
assign wn_re[1860] = 26'b00000000000000001101011010; assign wn_im[1860] = 26'b00000000000000001000101110; 
assign wn_re[1861] = 26'b00000000000000001101011100; assign wn_im[1861] = 26'b00000000000000001000101011; 
assign wn_re[1862] = 26'b00000000000000001101011101; assign wn_im[1862] = 26'b00000000000000001000101001; 
assign wn_re[1863] = 26'b00000000000000001101011111; assign wn_im[1863] = 26'b00000000000000001000100110; 
assign wn_re[1864] = 26'b00000000000000001101100001; assign wn_im[1864] = 26'b00000000000000001000100011; 
assign wn_re[1865] = 26'b00000000000000001101100010; assign wn_im[1865] = 26'b00000000000000001000100001; 
assign wn_re[1866] = 26'b00000000000000001101100100; assign wn_im[1866] = 26'b00000000000000001000011110; 
assign wn_re[1867] = 26'b00000000000000001101100110; assign wn_im[1867] = 26'b00000000000000001000011011; 
assign wn_re[1868] = 26'b00000000000000001101100111; assign wn_im[1868] = 26'b00000000000000001000011001; 
assign wn_re[1869] = 26'b00000000000000001101101001; assign wn_im[1869] = 26'b00000000000000001000010110; 
assign wn_re[1870] = 26'b00000000000000001101101011; assign wn_im[1870] = 26'b00000000000000001000010011; 
assign wn_re[1871] = 26'b00000000000000001101101100; assign wn_im[1871] = 26'b00000000000000001000010001; 
assign wn_re[1872] = 26'b00000000000000001101101110; assign wn_im[1872] = 26'b00000000000000001000001110; 
assign wn_re[1873] = 26'b00000000000000001101101111; assign wn_im[1873] = 26'b00000000000000001000001011; 
assign wn_re[1874] = 26'b00000000000000001101110001; assign wn_im[1874] = 26'b00000000000000001000001001; 
assign wn_re[1875] = 26'b00000000000000001101110011; assign wn_im[1875] = 26'b00000000000000001000000110; 
assign wn_re[1876] = 26'b00000000000000001101110100; assign wn_im[1876] = 26'b00000000000000001000000011; 
assign wn_re[1877] = 26'b00000000000000001101110110; assign wn_im[1877] = 26'b00000000000000001000000000; 
assign wn_re[1878] = 26'b00000000000000001101110111; assign wn_im[1878] = 26'b00000000000000000111111110; 
assign wn_re[1879] = 26'b00000000000000001101111001; assign wn_im[1879] = 26'b00000000000000000111111011; 
assign wn_re[1880] = 26'b00000000000000001101111010; assign wn_im[1880] = 26'b00000000000000000111111000; 
assign wn_re[1881] = 26'b00000000000000001101111100; assign wn_im[1881] = 26'b00000000000000000111110101; 
assign wn_re[1882] = 26'b00000000000000001101111110; assign wn_im[1882] = 26'b00000000000000000111110011; 
assign wn_re[1883] = 26'b00000000000000001101111111; assign wn_im[1883] = 26'b00000000000000000111110000; 
assign wn_re[1884] = 26'b00000000000000001110000001; assign wn_im[1884] = 26'b00000000000000000111101101; 
assign wn_re[1885] = 26'b00000000000000001110000010; assign wn_im[1885] = 26'b00000000000000000111101011; 
assign wn_re[1886] = 26'b00000000000000001110000100; assign wn_im[1886] = 26'b00000000000000000111101000; 
assign wn_re[1887] = 26'b00000000000000001110000101; assign wn_im[1887] = 26'b00000000000000000111100101; 
assign wn_re[1888] = 26'b00000000000000001110000111; assign wn_im[1888] = 26'b00000000000000000111100010; 
assign wn_re[1889] = 26'b00000000000000001110001000; assign wn_im[1889] = 26'b00000000000000000111011111; 
assign wn_re[1890] = 26'b00000000000000001110001010; assign wn_im[1890] = 26'b00000000000000000111011101; 
assign wn_re[1891] = 26'b00000000000000001110001011; assign wn_im[1891] = 26'b00000000000000000111011010; 
assign wn_re[1892] = 26'b00000000000000001110001100; assign wn_im[1892] = 26'b00000000000000000111010111; 
assign wn_re[1893] = 26'b00000000000000001110001110; assign wn_im[1893] = 26'b00000000000000000111010100; 
assign wn_re[1894] = 26'b00000000000000001110001111; assign wn_im[1894] = 26'b00000000000000000111010010; 
assign wn_re[1895] = 26'b00000000000000001110010001; assign wn_im[1895] = 26'b00000000000000000111001111; 
assign wn_re[1896] = 26'b00000000000000001110010010; assign wn_im[1896] = 26'b00000000000000000111001100; 
assign wn_re[1897] = 26'b00000000000000001110010100; assign wn_im[1897] = 26'b00000000000000000111001001; 
assign wn_re[1898] = 26'b00000000000000001110010101; assign wn_im[1898] = 26'b00000000000000000111000110; 
assign wn_re[1899] = 26'b00000000000000001110010110; assign wn_im[1899] = 26'b00000000000000000111000011; 
assign wn_re[1900] = 26'b00000000000000001110011000; assign wn_im[1900] = 26'b00000000000000000111000001; 
assign wn_re[1901] = 26'b00000000000000001110011001; assign wn_im[1901] = 26'b00000000000000000110111110; 
assign wn_re[1902] = 26'b00000000000000001110011010; assign wn_im[1902] = 26'b00000000000000000110111011; 
assign wn_re[1903] = 26'b00000000000000001110011100; assign wn_im[1903] = 26'b00000000000000000110111000; 
assign wn_re[1904] = 26'b00000000000000001110011101; assign wn_im[1904] = 26'b00000000000000000110110101; 
assign wn_re[1905] = 26'b00000000000000001110011111; assign wn_im[1905] = 26'b00000000000000000110110010; 
assign wn_re[1906] = 26'b00000000000000001110100000; assign wn_im[1906] = 26'b00000000000000000110110000; 
assign wn_re[1907] = 26'b00000000000000001110100001; assign wn_im[1907] = 26'b00000000000000000110101101; 
assign wn_re[1908] = 26'b00000000000000001110100010; assign wn_im[1908] = 26'b00000000000000000110101010; 
assign wn_re[1909] = 26'b00000000000000001110100100; assign wn_im[1909] = 26'b00000000000000000110100111; 
assign wn_re[1910] = 26'b00000000000000001110100101; assign wn_im[1910] = 26'b00000000000000000110100100; 
assign wn_re[1911] = 26'b00000000000000001110100110; assign wn_im[1911] = 26'b00000000000000000110100001; 
assign wn_re[1912] = 26'b00000000000000001110101000; assign wn_im[1912] = 26'b00000000000000000110011110; 
assign wn_re[1913] = 26'b00000000000000001110101001; assign wn_im[1913] = 26'b00000000000000000110011100; 
assign wn_re[1914] = 26'b00000000000000001110101010; assign wn_im[1914] = 26'b00000000000000000110011001; 
assign wn_re[1915] = 26'b00000000000000001110101011; assign wn_im[1915] = 26'b00000000000000000110010110; 
assign wn_re[1916] = 26'b00000000000000001110101101; assign wn_im[1916] = 26'b00000000000000000110010011; 
assign wn_re[1917] = 26'b00000000000000001110101110; assign wn_im[1917] = 26'b00000000000000000110010000; 
assign wn_re[1918] = 26'b00000000000000001110101111; assign wn_im[1918] = 26'b00000000000000000110001101; 
assign wn_re[1919] = 26'b00000000000000001110110000; assign wn_im[1919] = 26'b00000000000000000110001010; 
assign wn_re[1920] = 26'b00000000000000001110110010; assign wn_im[1920] = 26'b00000000000000000110000111; 
assign wn_re[1921] = 26'b00000000000000001110110011; assign wn_im[1921] = 26'b00000000000000000110000100; 
assign wn_re[1922] = 26'b00000000000000001110110100; assign wn_im[1922] = 26'b00000000000000000110000010; 
assign wn_re[1923] = 26'b00000000000000001110110101; assign wn_im[1923] = 26'b00000000000000000101111111; 
assign wn_re[1924] = 26'b00000000000000001110110110; assign wn_im[1924] = 26'b00000000000000000101111100; 
assign wn_re[1925] = 26'b00000000000000001110110111; assign wn_im[1925] = 26'b00000000000000000101111001; 
assign wn_re[1926] = 26'b00000000000000001110111001; assign wn_im[1926] = 26'b00000000000000000101110110; 
assign wn_re[1927] = 26'b00000000000000001110111010; assign wn_im[1927] = 26'b00000000000000000101110011; 
assign wn_re[1928] = 26'b00000000000000001110111011; assign wn_im[1928] = 26'b00000000000000000101110000; 
assign wn_re[1929] = 26'b00000000000000001110111100; assign wn_im[1929] = 26'b00000000000000000101101101; 
assign wn_re[1930] = 26'b00000000000000001110111101; assign wn_im[1930] = 26'b00000000000000000101101010; 
assign wn_re[1931] = 26'b00000000000000001110111110; assign wn_im[1931] = 26'b00000000000000000101100111; 
assign wn_re[1932] = 26'b00000000000000001110111111; assign wn_im[1932] = 26'b00000000000000000101100100; 
assign wn_re[1933] = 26'b00000000000000001111000000; assign wn_im[1933] = 26'b00000000000000000101100001; 
assign wn_re[1934] = 26'b00000000000000001111000010; assign wn_im[1934] = 26'b00000000000000000101011110; 
assign wn_re[1935] = 26'b00000000000000001111000011; assign wn_im[1935] = 26'b00000000000000000101011011; 
assign wn_re[1936] = 26'b00000000000000001111000100; assign wn_im[1936] = 26'b00000000000000000101011000; 
assign wn_re[1937] = 26'b00000000000000001111000101; assign wn_im[1937] = 26'b00000000000000000101010110; 
assign wn_re[1938] = 26'b00000000000000001111000110; assign wn_im[1938] = 26'b00000000000000000101010011; 
assign wn_re[1939] = 26'b00000000000000001111000111; assign wn_im[1939] = 26'b00000000000000000101010000; 
assign wn_re[1940] = 26'b00000000000000001111001000; assign wn_im[1940] = 26'b00000000000000000101001101; 
assign wn_re[1941] = 26'b00000000000000001111001001; assign wn_im[1941] = 26'b00000000000000000101001010; 
assign wn_re[1942] = 26'b00000000000000001111001010; assign wn_im[1942] = 26'b00000000000000000101000111; 
assign wn_re[1943] = 26'b00000000000000001111001011; assign wn_im[1943] = 26'b00000000000000000101000100; 
assign wn_re[1944] = 26'b00000000000000001111001100; assign wn_im[1944] = 26'b00000000000000000101000001; 
assign wn_re[1945] = 26'b00000000000000001111001101; assign wn_im[1945] = 26'b00000000000000000100111110; 
assign wn_re[1946] = 26'b00000000000000001111001110; assign wn_im[1946] = 26'b00000000000000000100111011; 
assign wn_re[1947] = 26'b00000000000000001111001111; assign wn_im[1947] = 26'b00000000000000000100111000; 
assign wn_re[1948] = 26'b00000000000000001111010000; assign wn_im[1948] = 26'b00000000000000000100110101; 
assign wn_re[1949] = 26'b00000000000000001111010001; assign wn_im[1949] = 26'b00000000000000000100110010; 
assign wn_re[1950] = 26'b00000000000000001111010010; assign wn_im[1950] = 26'b00000000000000000100101111; 
assign wn_re[1951] = 26'b00000000000000001111010010; assign wn_im[1951] = 26'b00000000000000000100101100; 
assign wn_re[1952] = 26'b00000000000000001111010011; assign wn_im[1952] = 26'b00000000000000000100101001; 
assign wn_re[1953] = 26'b00000000000000001111010100; assign wn_im[1953] = 26'b00000000000000000100100110; 
assign wn_re[1954] = 26'b00000000000000001111010101; assign wn_im[1954] = 26'b00000000000000000100100011; 
assign wn_re[1955] = 26'b00000000000000001111010110; assign wn_im[1955] = 26'b00000000000000000100100000; 
assign wn_re[1956] = 26'b00000000000000001111010111; assign wn_im[1956] = 26'b00000000000000000100011101; 
assign wn_re[1957] = 26'b00000000000000001111011000; assign wn_im[1957] = 26'b00000000000000000100011010; 
assign wn_re[1958] = 26'b00000000000000001111011001; assign wn_im[1958] = 26'b00000000000000000100010111; 
assign wn_re[1959] = 26'b00000000000000001111011010; assign wn_im[1959] = 26'b00000000000000000100010100; 
assign wn_re[1960] = 26'b00000000000000001111011010; assign wn_im[1960] = 26'b00000000000000000100010001; 
assign wn_re[1961] = 26'b00000000000000001111011011; assign wn_im[1961] = 26'b00000000000000000100001110; 
assign wn_re[1962] = 26'b00000000000000001111011100; assign wn_im[1962] = 26'b00000000000000000100001011; 
assign wn_re[1963] = 26'b00000000000000001111011101; assign wn_im[1963] = 26'b00000000000000000100001000; 
assign wn_re[1964] = 26'b00000000000000001111011110; assign wn_im[1964] = 26'b00000000000000000100000100; 
assign wn_re[1965] = 26'b00000000000000001111011110; assign wn_im[1965] = 26'b00000000000000000100000001; 
assign wn_re[1966] = 26'b00000000000000001111011111; assign wn_im[1966] = 26'b00000000000000000011111110; 
assign wn_re[1967] = 26'b00000000000000001111100000; assign wn_im[1967] = 26'b00000000000000000011111011; 
assign wn_re[1968] = 26'b00000000000000001111100001; assign wn_im[1968] = 26'b00000000000000000011111000; 
assign wn_re[1969] = 26'b00000000000000001111100010; assign wn_im[1969] = 26'b00000000000000000011110101; 
assign wn_re[1970] = 26'b00000000000000001111100010; assign wn_im[1970] = 26'b00000000000000000011110010; 
assign wn_re[1971] = 26'b00000000000000001111100011; assign wn_im[1971] = 26'b00000000000000000011101111; 
assign wn_re[1972] = 26'b00000000000000001111100100; assign wn_im[1972] = 26'b00000000000000000011101100; 
assign wn_re[1973] = 26'b00000000000000001111100101; assign wn_im[1973] = 26'b00000000000000000011101001; 
assign wn_re[1974] = 26'b00000000000000001111100101; assign wn_im[1974] = 26'b00000000000000000011100110; 
assign wn_re[1975] = 26'b00000000000000001111100110; assign wn_im[1975] = 26'b00000000000000000011100011; 
assign wn_re[1976] = 26'b00000000000000001111100111; assign wn_im[1976] = 26'b00000000000000000011100000; 
assign wn_re[1977] = 26'b00000000000000001111100111; assign wn_im[1977] = 26'b00000000000000000011011101; 
assign wn_re[1978] = 26'b00000000000000001111101000; assign wn_im[1978] = 26'b00000000000000000011011010; 
assign wn_re[1979] = 26'b00000000000000001111101001; assign wn_im[1979] = 26'b00000000000000000011010111; 
assign wn_re[1980] = 26'b00000000000000001111101001; assign wn_im[1980] = 26'b00000000000000000011010100; 
assign wn_re[1981] = 26'b00000000000000001111101010; assign wn_im[1981] = 26'b00000000000000000011010001; 
assign wn_re[1982] = 26'b00000000000000001111101011; assign wn_im[1982] = 26'b00000000000000000011001101; 
assign wn_re[1983] = 26'b00000000000000001111101011; assign wn_im[1983] = 26'b00000000000000000011001010; 
assign wn_re[1984] = 26'b00000000000000001111101100; assign wn_im[1984] = 26'b00000000000000000011000111; 
assign wn_re[1985] = 26'b00000000000000001111101100; assign wn_im[1985] = 26'b00000000000000000011000100; 
assign wn_re[1986] = 26'b00000000000000001111101101; assign wn_im[1986] = 26'b00000000000000000011000001; 
assign wn_re[1987] = 26'b00000000000000001111101110; assign wn_im[1987] = 26'b00000000000000000010111110; 
assign wn_re[1988] = 26'b00000000000000001111101110; assign wn_im[1988] = 26'b00000000000000000010111011; 
assign wn_re[1989] = 26'b00000000000000001111101111; assign wn_im[1989] = 26'b00000000000000000010111000; 
assign wn_re[1990] = 26'b00000000000000001111101111; assign wn_im[1990] = 26'b00000000000000000010110101; 
assign wn_re[1991] = 26'b00000000000000001111110000; assign wn_im[1991] = 26'b00000000000000000010110010; 
assign wn_re[1992] = 26'b00000000000000001111110000; assign wn_im[1992] = 26'b00000000000000000010101111; 
assign wn_re[1993] = 26'b00000000000000001111110001; assign wn_im[1993] = 26'b00000000000000000010101011; 
assign wn_re[1994] = 26'b00000000000000001111110001; assign wn_im[1994] = 26'b00000000000000000010101000; 
assign wn_re[1995] = 26'b00000000000000001111110010; assign wn_im[1995] = 26'b00000000000000000010100101; 
assign wn_re[1996] = 26'b00000000000000001111110010; assign wn_im[1996] = 26'b00000000000000000010100010; 
assign wn_re[1997] = 26'b00000000000000001111110011; assign wn_im[1997] = 26'b00000000000000000010011111; 
assign wn_re[1998] = 26'b00000000000000001111110011; assign wn_im[1998] = 26'b00000000000000000010011100; 
assign wn_re[1999] = 26'b00000000000000001111110100; assign wn_im[1999] = 26'b00000000000000000010011001; 
assign wn_re[2000] = 26'b00000000000000001111110100; assign wn_im[2000] = 26'b00000000000000000010010110; 
assign wn_re[2001] = 26'b00000000000000001111110101; assign wn_im[2001] = 26'b00000000000000000010010011; 
assign wn_re[2002] = 26'b00000000000000001111110101; assign wn_im[2002] = 26'b00000000000000000010010000; 
assign wn_re[2003] = 26'b00000000000000001111110110; assign wn_im[2003] = 26'b00000000000000000010001100; 
assign wn_re[2004] = 26'b00000000000000001111110110; assign wn_im[2004] = 26'b00000000000000000010001001; 
assign wn_re[2005] = 26'b00000000000000001111110111; assign wn_im[2005] = 26'b00000000000000000010000110; 
assign wn_re[2006] = 26'b00000000000000001111110111; assign wn_im[2006] = 26'b00000000000000000010000011; 
assign wn_re[2007] = 26'b00000000000000001111110111; assign wn_im[2007] = 26'b00000000000000000010000000; 
assign wn_re[2008] = 26'b00000000000000001111111000; assign wn_im[2008] = 26'b00000000000000000001111101; 
assign wn_re[2009] = 26'b00000000000000001111111000; assign wn_im[2009] = 26'b00000000000000000001111010; 
assign wn_re[2010] = 26'b00000000000000001111111001; assign wn_im[2010] = 26'b00000000000000000001110111; 
assign wn_re[2011] = 26'b00000000000000001111111001; assign wn_im[2011] = 26'b00000000000000000001110011; 
assign wn_re[2012] = 26'b00000000000000001111111001; assign wn_im[2012] = 26'b00000000000000000001110000; 
assign wn_re[2013] = 26'b00000000000000001111111010; assign wn_im[2013] = 26'b00000000000000000001101101; 
assign wn_re[2014] = 26'b00000000000000001111111010; assign wn_im[2014] = 26'b00000000000000000001101010; 
assign wn_re[2015] = 26'b00000000000000001111111010; assign wn_im[2015] = 26'b00000000000000000001100111; 
assign wn_re[2016] = 26'b00000000000000001111111011; assign wn_im[2016] = 26'b00000000000000000001100100; 
assign wn_re[2017] = 26'b00000000000000001111111011; assign wn_im[2017] = 26'b00000000000000000001100001; 
assign wn_re[2018] = 26'b00000000000000001111111011; assign wn_im[2018] = 26'b00000000000000000001011110; 
assign wn_re[2019] = 26'b00000000000000001111111011; assign wn_im[2019] = 26'b00000000000000000001011010; 
assign wn_re[2020] = 26'b00000000000000001111111100; assign wn_im[2020] = 26'b00000000000000000001010111; 
assign wn_re[2021] = 26'b00000000000000001111111100; assign wn_im[2021] = 26'b00000000000000000001010100; 
assign wn_re[2022] = 26'b00000000000000001111111100; assign wn_im[2022] = 26'b00000000000000000001010001; 
assign wn_re[2023] = 26'b00000000000000001111111100; assign wn_im[2023] = 26'b00000000000000000001001110; 
assign wn_re[2024] = 26'b00000000000000001111111101; assign wn_im[2024] = 26'b00000000000000000001001011; 
assign wn_re[2025] = 26'b00000000000000001111111101; assign wn_im[2025] = 26'b00000000000000000001001000; 
assign wn_re[2026] = 26'b00000000000000001111111101; assign wn_im[2026] = 26'b00000000000000000001000101; 
assign wn_re[2027] = 26'b00000000000000001111111101; assign wn_im[2027] = 26'b00000000000000000001000001; 
assign wn_re[2028] = 26'b00000000000000001111111110; assign wn_im[2028] = 26'b00000000000000000000111110; 
assign wn_re[2029] = 26'b00000000000000001111111110; assign wn_im[2029] = 26'b00000000000000000000111011; 
assign wn_re[2030] = 26'b00000000000000001111111110; assign wn_im[2030] = 26'b00000000000000000000111000; 
assign wn_re[2031] = 26'b00000000000000001111111110; assign wn_im[2031] = 26'b00000000000000000000110101; 
assign wn_re[2032] = 26'b00000000000000001111111110; assign wn_im[2032] = 26'b00000000000000000000110010; 
assign wn_re[2033] = 26'b00000000000000001111111110; assign wn_im[2033] = 26'b00000000000000000000101111; 
assign wn_re[2034] = 26'b00000000000000001111111111; assign wn_im[2034] = 26'b00000000000000000000101011; 
assign wn_re[2035] = 26'b00000000000000001111111111; assign wn_im[2035] = 26'b00000000000000000000101000; 
assign wn_re[2036] = 26'b00000000000000001111111111; assign wn_im[2036] = 26'b00000000000000000000100101; 
assign wn_re[2037] = 26'b00000000000000001111111111; assign wn_im[2037] = 26'b00000000000000000000100010; 
assign wn_re[2038] = 26'b00000000000000001111111111; assign wn_im[2038] = 26'b00000000000000000000011111; 
assign wn_re[2039] = 26'b00000000000000001111111111; assign wn_im[2039] = 26'b00000000000000000000011100; 
assign wn_re[2040] = 26'b00000000000000001111111111; assign wn_im[2040] = 26'b00000000000000000000011001; 
assign wn_re[2041] = 26'b00000000000000001111111111; assign wn_im[2041] = 26'b00000000000000000000010101; 
assign wn_re[2042] = 26'b00000000000000001111111111; assign wn_im[2042] = 26'b00000000000000000000010010; 
assign wn_re[2043] = 26'b00000000000000001111111111; assign wn_im[2043] = 26'b00000000000000000000001111; 
assign wn_re[2044] = 26'b00000000000000001111111111; assign wn_im[2044] = 26'b00000000000000000000001100; 
assign wn_re[2045] = 26'b00000000000000001111111111; assign wn_im[2045] = 26'b00000000000000000000001001; 
assign wn_re[2046] = 26'b00000000000000001111111111; assign wn_im[2046] = 26'b00000000000000000000000110; 
assign wn_re[2047] = 26'b00000000000000001111111111; assign wn_im[2047] = 26'b00000000000000000000000011; 

endmodule
