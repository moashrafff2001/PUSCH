module phi4 (
        input   [4:0]   u,   //  Sequence number
        input   [9:0]   counter,   //  Counter of the generator
        output  [1:0]  phi_value  //  phase of the sequence
    );

    wire [1:0] phi4 [0:29][0:23];
    assign phi_value = phi4[u][counter];
assign phi4 [0][0] = 2'b10;
assign phi4 [0][1] = 2'b11;
assign phi4 [0][2] = 2'b01;
assign phi4 [0][3] = 2'b10;
assign phi4 [0][4] = 2'b01;
assign phi4 [0][5] = 2'b00;
assign phi4 [0][6] = 2'b01;
assign phi4 [0][7] = 2'b10;
assign phi4 [0][8] = 2'b00;
assign phi4 [0][9] = 2'b11;
assign phi4 [0][10] = 2'b10;
assign phi4 [0][11] = 2'b11;
assign phi4 [0][12] = 2'b10;
assign phi4 [0][13] = 2'b00;
assign phi4 [0][14] = 2'b01;
assign phi4 [0][15] = 2'b11;
assign phi4 [0][16] = 2'b10;
assign phi4 [0][17] = 2'b11;
assign phi4 [0][18] = 2'b01;
assign phi4 [0][19] = 2'b01;
assign phi4 [0][20] = 2'b01;
assign phi4 [0][21] = 2'b11;
assign phi4 [0][22] = 2'b11;
assign phi4 [0][23] = 2'b11;
assign phi4 [1][0] = 2'b10;
assign phi4 [1][1] = 2'b11;
assign phi4 [1][2] = 2'b01;
assign phi4 [1][3] = 2'b00;
assign phi4 [1][4] = 2'b00;
assign phi4 [1][5] = 2'b11;
assign phi4 [1][6] = 2'b00;
assign phi4 [1][7] = 2'b11;
assign phi4 [1][8] = 2'b11;
assign phi4 [1][9] = 2'b00;
assign phi4 [1][10] = 2'b11;
assign phi4 [1][11] = 2'b10;
assign phi4 [1][12] = 2'b10;
assign phi4 [1][13] = 2'b01;
assign phi4 [1][14] = 2'b11;
assign phi4 [1][15] = 2'b01;
assign phi4 [1][16] = 2'b01;
assign phi4 [1][17] = 2'b01;
assign phi4 [1][18] = 2'b11;
assign phi4 [1][19] = 2'b00;
assign phi4 [1][20] = 2'b01;
assign phi4 [1][21] = 2'b01;
assign phi4 [1][22] = 2'b11;
assign phi4 [1][23] = 2'b11;
assign phi4 [2][0] = 2'b10;
assign phi4 [2][1] = 2'b11;
assign phi4 [2][2] = 2'b11;
assign phi4 [2][3] = 2'b00;
assign phi4 [2][4] = 2'b10;
assign phi4 [2][5] = 2'b10;
assign phi4 [2][6] = 2'b11;
assign phi4 [2][7] = 2'b00;
assign phi4 [2][8] = 2'b01;
assign phi4 [2][9] = 2'b10;
assign phi4 [2][10] = 2'b11;
assign phi4 [2][11] = 2'b10;
assign phi4 [2][12] = 2'b10;
assign phi4 [2][13] = 2'b11;
assign phi4 [2][14] = 2'b00;
assign phi4 [2][15] = 2'b00;
assign phi4 [2][16] = 2'b01;
assign phi4 [2][17] = 2'b00;
assign phi4 [2][18] = 2'b11;
assign phi4 [2][19] = 2'b10;
assign phi4 [2][20] = 2'b10;
assign phi4 [2][21] = 2'b01;
assign phi4 [2][22] = 2'b11;
assign phi4 [2][23] = 2'b11;
assign phi4 [3][0] = 2'b00;
assign phi4 [3][1] = 2'b11;
assign phi4 [3][2] = 2'b01;
assign phi4 [3][3] = 2'b10;
assign phi4 [3][4] = 2'b11;
assign phi4 [3][5] = 2'b10;
assign phi4 [3][6] = 2'b01;
assign phi4 [3][7] = 2'b01;
assign phi4 [3][8] = 2'b00;
assign phi4 [3][9] = 2'b10;
assign phi4 [3][10] = 2'b00;
assign phi4 [3][11] = 2'b00;
assign phi4 [3][12] = 2'b01;
assign phi4 [3][13] = 2'b11;
assign phi4 [3][14] = 2'b10;
assign phi4 [3][15] = 2'b11;
assign phi4 [3][16] = 2'b11;
assign phi4 [3][17] = 2'b11;
assign phi4 [3][18] = 2'b10;
assign phi4 [3][19] = 2'b01;
assign phi4 [3][20] = 2'b11;
assign phi4 [3][21] = 2'b10;
assign phi4 [3][22] = 2'b11;
assign phi4 [3][23] = 2'b11;
assign phi4 [4][0] = 2'b10;
assign phi4 [4][1] = 2'b01;
assign phi4 [4][2] = 2'b11;
assign phi4 [4][3] = 2'b11;
assign phi4 [4][4] = 2'b10;
assign phi4 [4][5] = 2'b01;
assign phi4 [4][6] = 2'b10;
assign phi4 [4][7] = 2'b10;
assign phi4 [4][8] = 2'b00;
assign phi4 [4][9] = 2'b01;
assign phi4 [4][10] = 2'b00;
assign phi4 [4][11] = 2'b01;
assign phi4 [4][12] = 2'b10;
assign phi4 [4][13] = 2'b10;
assign phi4 [4][14] = 2'b11;
assign phi4 [4][15] = 2'b00;
assign phi4 [4][16] = 2'b01;
assign phi4 [4][17] = 2'b00;
assign phi4 [4][18] = 2'b10;
assign phi4 [4][19] = 2'b11;
assign phi4 [4][20] = 2'b00;
assign phi4 [4][21] = 2'b10;
assign phi4 [4][22] = 2'b11;
assign phi4 [4][23] = 2'b11;
assign phi4 [5][0] = 2'b11;
assign phi4 [5][1] = 2'b10;
assign phi4 [5][2] = 2'b00;
assign phi4 [5][3] = 2'b11;
assign phi4 [5][4] = 2'b11;
assign phi4 [5][5] = 2'b00;
assign phi4 [5][6] = 2'b00;
assign phi4 [5][7] = 2'b11;
assign phi4 [5][8] = 2'b01;
assign phi4 [5][9] = 2'b10;
assign phi4 [5][10] = 2'b10;
assign phi4 [5][11] = 2'b11;
assign phi4 [5][12] = 2'b00;
assign phi4 [5][13] = 2'b01;
assign phi4 [5][14] = 2'b00;
assign phi4 [5][15] = 2'b10;
assign phi4 [5][16] = 2'b11;
assign phi4 [5][17] = 2'b10;
assign phi4 [5][18] = 2'b11;
assign phi4 [5][19] = 2'b00;
assign phi4 [5][20] = 2'b11;
assign phi4 [5][21] = 2'b11;
assign phi4 [5][22] = 2'b11;
assign phi4 [5][23] = 2'b11;
assign phi4 [6][0] = 2'b11;
assign phi4 [6][1] = 2'b01;
assign phi4 [6][2] = 2'b00;
assign phi4 [6][3] = 2'b01;
assign phi4 [6][4] = 2'b10;
assign phi4 [6][5] = 2'b00;
assign phi4 [6][6] = 2'b11;
assign phi4 [6][7] = 2'b00;
assign phi4 [6][8] = 2'b11;
assign phi4 [6][9] = 2'b00;
assign phi4 [6][10] = 2'b10;
assign phi4 [6][11] = 2'b11;
assign phi4 [6][12] = 2'b10;
assign phi4 [6][13] = 2'b11;
assign phi4 [6][14] = 2'b11;
assign phi4 [6][15] = 2'b11;
assign phi4 [6][16] = 2'b11;
assign phi4 [6][17] = 2'b10;
assign phi4 [6][18] = 2'b10;
assign phi4 [6][19] = 2'b10;
assign phi4 [6][20] = 2'b00;
assign phi4 [6][21] = 2'b00;
assign phi4 [6][22] = 2'b11;
assign phi4 [6][23] = 2'b11;
assign phi4 [7][0] = 2'b11;
assign phi4 [7][1] = 2'b00;
assign phi4 [7][2] = 2'b01;
assign phi4 [7][3] = 2'b10;
assign phi4 [7][4] = 2'b00;
assign phi4 [7][5] = 2'b10;
assign phi4 [7][6] = 2'b01;
assign phi4 [7][7] = 2'b11;
assign phi4 [7][8] = 2'b01;
assign phi4 [7][9] = 2'b10;
assign phi4 [7][10] = 2'b11;
assign phi4 [7][11] = 2'b10;
assign phi4 [7][12] = 2'b11;
assign phi4 [7][13] = 2'b01;
assign phi4 [7][14] = 2'b10;
assign phi4 [7][15] = 2'b10;
assign phi4 [7][16] = 2'b10;
assign phi4 [7][17] = 2'b11;
assign phi4 [7][18] = 2'b10;
assign phi4 [7][19] = 2'b10;
assign phi4 [7][20] = 2'b11;
assign phi4 [7][21] = 2'b01;
assign phi4 [7][22] = 2'b01;
assign phi4 [7][23] = 2'b11;
assign phi4 [8][0] = 2'b11;
assign phi4 [8][1] = 2'b00;
assign phi4 [8][2] = 2'b11;
assign phi4 [8][3] = 2'b01;
assign phi4 [8][4] = 2'b10;
assign phi4 [8][5] = 2'b10;
assign phi4 [8][6] = 2'b10;
assign phi4 [8][7] = 2'b11;
assign phi4 [8][8] = 2'b01;
assign phi4 [8][9] = 2'b00;
assign phi4 [8][10] = 2'b10;
assign phi4 [8][11] = 2'b11;
assign phi4 [8][12] = 2'b10;
assign phi4 [8][13] = 2'b00;
assign phi4 [8][14] = 2'b01;
assign phi4 [8][15] = 2'b10;
assign phi4 [8][16] = 2'b00;
assign phi4 [8][17] = 2'b10;
assign phi4 [8][18] = 2'b00;
assign phi4 [8][19] = 2'b11;
assign phi4 [8][20] = 2'b11;
assign phi4 [8][21] = 2'b11;
assign phi4 [8][22] = 2'b11;
assign phi4 [8][23] = 2'b11;
assign phi4 [9][0] = 2'b00;
assign phi4 [9][1] = 2'b00;
assign phi4 [9][2] = 2'b10;
assign phi4 [9][3] = 2'b11;
assign phi4 [9][4] = 2'b10;
assign phi4 [9][5] = 2'b00;
assign phi4 [9][6] = 2'b00;
assign phi4 [9][7] = 2'b11;
assign phi4 [9][8] = 2'b00;
assign phi4 [9][9] = 2'b10;
assign phi4 [9][10] = 2'b00;
assign phi4 [9][11] = 2'b11;
assign phi4 [9][12] = 2'b01;
assign phi4 [9][13] = 2'b11;
assign phi4 [9][14] = 2'b11;
assign phi4 [9][15] = 2'b01;
assign phi4 [9][16] = 2'b10;
assign phi4 [9][17] = 2'b11;
assign phi4 [9][18] = 2'b00;
assign phi4 [9][19] = 2'b01;
assign phi4 [9][20] = 2'b11;
assign phi4 [9][21] = 2'b00;
assign phi4 [9][22] = 2'b11;
assign phi4 [9][23] = 2'b11;
assign phi4 [10][0] = 2'b11;
assign phi4 [10][1] = 2'b11;
assign phi4 [10][2] = 2'b11;
assign phi4 [10][3] = 2'b10;
assign phi4 [10][4] = 2'b01;
assign phi4 [10][5] = 2'b11;
assign phi4 [10][6] = 2'b01;
assign phi4 [10][7] = 2'b00;
assign phi4 [10][8] = 2'b01;
assign phi4 [10][9] = 2'b00;
assign phi4 [10][10] = 2'b11;
assign phi4 [10][11] = 2'b10;
assign phi4 [10][12] = 2'b10;
assign phi4 [10][13] = 2'b11;
assign phi4 [10][14] = 2'b00;
assign phi4 [10][15] = 2'b00;
assign phi4 [10][16] = 2'b01;
assign phi4 [10][17] = 2'b00;
assign phi4 [10][18] = 2'b10;
assign phi4 [10][19] = 2'b11;
assign phi4 [10][20] = 2'b01;
assign phi4 [10][21] = 2'b00;
assign phi4 [10][22] = 2'b01;
assign phi4 [10][23] = 2'b11;
assign phi4 [11][0] = 2'b11;
assign phi4 [11][1] = 2'b01;
assign phi4 [11][2] = 2'b10;
assign phi4 [11][3] = 2'b01;
assign phi4 [11][4] = 2'b00;
assign phi4 [11][5] = 2'b10;
assign phi4 [11][6] = 2'b10;
assign phi4 [11][7] = 2'b10;
assign phi4 [11][8] = 2'b01;
assign phi4 [11][9] = 2'b01;
assign phi4 [11][10] = 2'b00;
assign phi4 [11][11] = 2'b00;
assign phi4 [11][12] = 2'b00;
assign phi4 [11][13] = 2'b01;
assign phi4 [11][14] = 2'b01;
assign phi4 [11][15] = 2'b00;
assign phi4 [11][16] = 2'b11;
assign phi4 [11][17] = 2'b11;
assign phi4 [11][18] = 2'b10;
assign phi4 [11][19] = 2'b00;
assign phi4 [11][20] = 2'b11;
assign phi4 [11][21] = 2'b00;
assign phi4 [11][22] = 2'b01;
assign phi4 [11][23] = 2'b11;
assign phi4 [12][0] = 2'b01;
assign phi4 [12][1] = 2'b11;
assign phi4 [12][2] = 2'b01;
assign phi4 [12][3] = 2'b10;
assign phi4 [12][4] = 2'b11;
assign phi4 [12][5] = 2'b00;
assign phi4 [12][6] = 2'b01;
assign phi4 [12][7] = 2'b00;
assign phi4 [12][8] = 2'b10;
assign phi4 [12][9] = 2'b10;
assign phi4 [12][10] = 2'b11;
assign phi4 [12][11] = 2'b10;
assign phi4 [12][12] = 2'b01;
assign phi4 [12][13] = 2'b11;
assign phi4 [12][14] = 2'b01;
assign phi4 [12][15] = 2'b10;
assign phi4 [12][16] = 2'b10;
assign phi4 [12][17] = 2'b01;
assign phi4 [12][18] = 2'b01;
assign phi4 [12][19] = 2'b11;
assign phi4 [12][20] = 2'b11;
assign phi4 [12][21] = 2'b01;
assign phi4 [12][22] = 2'b11;
assign phi4 [12][23] = 2'b11;
assign phi4 [13][0] = 2'b11;
assign phi4 [13][1] = 2'b01;
assign phi4 [13][2] = 2'b10;
assign phi4 [13][3] = 2'b01;
assign phi4 [13][4] = 2'b10;
assign phi4 [13][5] = 2'b01;
assign phi4 [13][6] = 2'b01;
assign phi4 [13][7] = 2'b00;
assign phi4 [13][8] = 2'b00;
assign phi4 [13][9] = 2'b11;
assign phi4 [13][10] = 2'b00;
assign phi4 [13][11] = 2'b01;
assign phi4 [13][12] = 2'b11;
assign phi4 [13][13] = 2'b01;
assign phi4 [13][14] = 2'b11;
assign phi4 [13][15] = 2'b11;
assign phi4 [13][16] = 2'b10;
assign phi4 [13][17] = 2'b00;
assign phi4 [13][18] = 2'b01;
assign phi4 [13][19] = 2'b11;
assign phi4 [13][20] = 2'b10;
assign phi4 [13][21] = 2'b10;
assign phi4 [13][22] = 2'b11;
assign phi4 [13][23] = 2'b11;
assign phi4 [14][0] = 2'b11;
assign phi4 [14][1] = 2'b00;
assign phi4 [14][2] = 2'b11;
assign phi4 [14][3] = 2'b10;
assign phi4 [14][4] = 2'b10;
assign phi4 [14][5] = 2'b01;
assign phi4 [14][6] = 2'b00;
assign phi4 [14][7] = 2'b01;
assign phi4 [14][8] = 2'b11;
assign phi4 [14][9] = 2'b00;
assign phi4 [14][10] = 2'b10;
assign phi4 [14][11] = 2'b01;
assign phi4 [14][12] = 2'b01;
assign phi4 [14][13] = 2'b10;
assign phi4 [14][14] = 2'b11;
assign phi4 [14][15] = 2'b01;
assign phi4 [14][16] = 2'b11;
assign phi4 [14][17] = 2'b10;
assign phi4 [14][18] = 2'b10;
assign phi4 [14][19] = 2'b11;
assign phi4 [14][20] = 2'b11;
assign phi4 [14][21] = 2'b11;
assign phi4 [14][22] = 2'b01;
assign phi4 [14][23] = 2'b11;
assign phi4 [15][0] = 2'b11;
assign phi4 [15][1] = 2'b10;
assign phi4 [15][2] = 2'b10;
assign phi4 [15][3] = 2'b11;
assign phi4 [15][4] = 2'b00;
assign phi4 [15][5] = 2'b11;
assign phi4 [15][6] = 2'b11;
assign phi4 [15][7] = 2'b10;
assign phi4 [15][8] = 2'b10;
assign phi4 [15][9] = 2'b01;
assign phi4 [15][10] = 2'b10;
assign phi4 [15][11] = 2'b00;
assign phi4 [15][12] = 2'b10;
assign phi4 [15][13] = 2'b01;
assign phi4 [15][14] = 2'b00;
assign phi4 [15][15] = 2'b11;
assign phi4 [15][16] = 2'b10;
assign phi4 [15][17] = 2'b01;
assign phi4 [15][18] = 2'b00;
assign phi4 [15][19] = 2'b00;
assign phi4 [15][20] = 2'b10;
assign phi4 [15][21] = 2'b10;
assign phi4 [15][22] = 2'b11;
assign phi4 [15][23] = 2'b11;
assign phi4 [16][0] = 2'b11;
assign phi4 [16][1] = 2'b11;
assign phi4 [16][2] = 2'b00;
assign phi4 [16][3] = 2'b10;
assign phi4 [16][4] = 2'b01;
assign phi4 [16][5] = 2'b01;
assign phi4 [16][6] = 2'b11;
assign phi4 [16][7] = 2'b10;
assign phi4 [16][8] = 2'b00;
assign phi4 [16][9] = 2'b10;
assign phi4 [16][10] = 2'b10;
assign phi4 [16][11] = 2'b00;
assign phi4 [16][12] = 2'b00;
assign phi4 [16][13] = 2'b10;
assign phi4 [16][14] = 2'b10;
assign phi4 [16][15] = 2'b01;
assign phi4 [16][16] = 2'b11;
assign phi4 [16][17] = 2'b00;
assign phi4 [16][18] = 2'b11;
assign phi4 [16][19] = 2'b00;
assign phi4 [16][20] = 2'b10;
assign phi4 [16][21] = 2'b10;
assign phi4 [16][22] = 2'b10;
assign phi4 [16][23] = 2'b11;
assign phi4 [17][0] = 2'b01;
assign phi4 [17][1] = 2'b10;
assign phi4 [17][2] = 2'b01;
assign phi4 [17][3] = 2'b10;
assign phi4 [17][4] = 2'b00;
assign phi4 [17][5] = 2'b11;
assign phi4 [17][6] = 2'b00;
assign phi4 [17][7] = 2'b00;
assign phi4 [17][8] = 2'b11;
assign phi4 [17][9] = 2'b11;
assign phi4 [17][10] = 2'b01;
assign phi4 [17][11] = 2'b11;
assign phi4 [17][12] = 2'b10;
assign phi4 [17][13] = 2'b10;
assign phi4 [17][14] = 2'b10;
assign phi4 [17][15] = 2'b10;
assign phi4 [17][16] = 2'b10;
assign phi4 [17][17] = 2'b11;
assign phi4 [17][18] = 2'b11;
assign phi4 [17][19] = 2'b10;
assign phi4 [17][20] = 2'b00;
assign phi4 [17][21] = 2'b00;
assign phi4 [17][22] = 2'b11;
assign phi4 [17][23] = 2'b11;
assign phi4 [18][0] = 2'b11;
assign phi4 [18][1] = 2'b00;
assign phi4 [18][2] = 2'b11;
assign phi4 [18][3] = 2'b00;
assign phi4 [18][4] = 2'b11;
assign phi4 [18][5] = 2'b11;
assign phi4 [18][6] = 2'b00;
assign phi4 [18][7] = 2'b11;
assign phi4 [18][8] = 2'b00;
assign phi4 [18][9] = 2'b11;
assign phi4 [18][10] = 2'b11;
assign phi4 [18][11] = 2'b11;
assign phi4 [18][12] = 2'b11;
assign phi4 [18][13] = 2'b11;
assign phi4 [18][14] = 2'b00;
assign phi4 [18][15] = 2'b11;
assign phi4 [18][16] = 2'b11;
assign phi4 [18][17] = 2'b00;
assign phi4 [18][18] = 2'b00;
assign phi4 [18][19] = 2'b11;
assign phi4 [18][20] = 2'b00;
assign phi4 [18][21] = 2'b00;
assign phi4 [18][22] = 2'b11;
assign phi4 [18][23] = 2'b11;
assign phi4 [19][0] = 2'b11;
assign phi4 [19][1] = 2'b11;
assign phi4 [19][2] = 2'b01;
assign phi4 [19][3] = 2'b01;
assign phi4 [19][4] = 2'b00;
assign phi4 [19][5] = 2'b10;
assign phi4 [19][6] = 2'b10;
assign phi4 [19][7] = 2'b10;
assign phi4 [19][8] = 2'b00;
assign phi4 [19][9] = 2'b11;
assign phi4 [19][10] = 2'b10;
assign phi4 [19][11] = 2'b00;
assign phi4 [19][12] = 2'b10;
assign phi4 [19][13] = 2'b01;
assign phi4 [19][14] = 2'b11;
assign phi4 [19][15] = 2'b10;
assign phi4 [19][16] = 2'b11;
assign phi4 [19][17] = 2'b10;
assign phi4 [19][18] = 2'b10;
assign phi4 [19][19] = 2'b00;
assign phi4 [19][20] = 2'b11;
assign phi4 [19][21] = 2'b01;
assign phi4 [19][22] = 2'b10;
assign phi4 [19][23] = 2'b11;
assign phi4 [20][0] = 2'b11;
assign phi4 [20][1] = 2'b11;
assign phi4 [20][2] = 2'b10;
assign phi4 [20][3] = 2'b10;
assign phi4 [20][4] = 2'b10;
assign phi4 [20][5] = 2'b11;
assign phi4 [20][6] = 2'b00;
assign phi4 [20][7] = 2'b10;
assign phi4 [20][8] = 2'b11;
assign phi4 [20][9] = 2'b10;
assign phi4 [20][10] = 2'b01;
assign phi4 [20][11] = 2'b11;
assign phi4 [20][12] = 2'b00;
assign phi4 [20][13] = 2'b11;
assign phi4 [20][14] = 2'b01;
assign phi4 [20][15] = 2'b11;
assign phi4 [20][16] = 2'b01;
assign phi4 [20][17] = 2'b01;
assign phi4 [20][18] = 2'b00;
assign phi4 [20][19] = 2'b10;
assign phi4 [20][20] = 2'b10;
assign phi4 [20][21] = 2'b00;
assign phi4 [20][22] = 2'b11;
assign phi4 [20][23] = 2'b11;
assign phi4 [21][0] = 2'b01;
assign phi4 [21][1] = 2'b10;
assign phi4 [21][2] = 2'b00;
assign phi4 [21][3] = 2'b10;
assign phi4 [21][4] = 2'b01;
assign phi4 [21][5] = 2'b11;
assign phi4 [21][6] = 2'b00;
assign phi4 [21][7] = 2'b00;
assign phi4 [21][8] = 2'b01;
assign phi4 [21][9] = 2'b10;
assign phi4 [21][10] = 2'b11;
assign phi4 [21][11] = 2'b01;
assign phi4 [21][12] = 2'b00;
assign phi4 [21][13] = 2'b11;
assign phi4 [21][14] = 2'b01;
assign phi4 [21][15] = 2'b10;
assign phi4 [21][16] = 2'b10;
assign phi4 [21][17] = 2'b10;
assign phi4 [21][18] = 2'b10;
assign phi4 [21][19] = 2'b00;
assign phi4 [21][20] = 2'b11;
assign phi4 [21][21] = 2'b11;
assign phi4 [21][22] = 2'b11;
assign phi4 [21][23] = 2'b11;
assign phi4 [22][0] = 2'b11;
assign phi4 [22][1] = 2'b00;
assign phi4 [22][2] = 2'b11;
assign phi4 [22][3] = 2'b01;
assign phi4 [22][4] = 2'b11;
assign phi4 [22][5] = 2'b00;
assign phi4 [22][6] = 2'b11;
assign phi4 [22][7] = 2'b01;
assign phi4 [22][8] = 2'b00;
assign phi4 [22][9] = 2'b10;
assign phi4 [22][10] = 2'b11;
assign phi4 [22][11] = 2'b10;
assign phi4 [22][12] = 2'b11;
assign phi4 [22][13] = 2'b11;
assign phi4 [22][14] = 2'b11;
assign phi4 [22][15] = 2'b11;
assign phi4 [22][16] = 2'b00;
assign phi4 [22][17] = 2'b01;
assign phi4 [22][18] = 2'b10;
assign phi4 [22][19] = 2'b00;
assign phi4 [22][20] = 2'b01;
assign phi4 [22][21] = 2'b01;
assign phi4 [22][22] = 2'b01;
assign phi4 [22][23] = 2'b11;
assign phi4 [23][0] = 2'b11;
assign phi4 [23][1] = 2'b10;
assign phi4 [23][2] = 2'b00;
assign phi4 [23][3] = 2'b11;
assign phi4 [23][4] = 2'b10;
assign phi4 [23][5] = 2'b10;
assign phi4 [23][6] = 2'b00;
assign phi4 [23][7] = 2'b00;
assign phi4 [23][8] = 2'b00;
assign phi4 [23][9] = 2'b01;
assign phi4 [23][10] = 2'b01;
assign phi4 [23][11] = 2'b10;
assign phi4 [23][12] = 2'b00;
assign phi4 [23][13] = 2'b10;
assign phi4 [23][14] = 2'b00;
assign phi4 [23][15] = 2'b10;
assign phi4 [23][16] = 2'b10;
assign phi4 [23][17] = 2'b11;
assign phi4 [23][18] = 2'b11;
assign phi4 [23][19] = 2'b11;
assign phi4 [23][20] = 2'b01;
assign phi4 [23][21] = 2'b00;
assign phi4 [23][22] = 2'b10;
assign phi4 [23][23] = 2'b11;
assign phi4 [24][0] = 2'b11;
assign phi4 [24][1] = 2'b01;
assign phi4 [24][2] = 2'b10;
assign phi4 [24][3] = 2'b11;
assign phi4 [24][4] = 2'b10;
assign phi4 [24][5] = 2'b10;
assign phi4 [24][6] = 2'b10;
assign phi4 [24][7] = 2'b01;
assign phi4 [24][8] = 2'b10;
assign phi4 [24][9] = 2'b10;
assign phi4 [24][10] = 2'b01;
assign phi4 [24][11] = 2'b11;
assign phi4 [24][12] = 2'b10;
assign phi4 [24][13] = 2'b01;
assign phi4 [24][14] = 2'b11;
assign phi4 [24][15] = 2'b01;
assign phi4 [24][16] = 2'b11;
assign phi4 [24][17] = 2'b10;
assign phi4 [24][18] = 2'b01;
assign phi4 [24][19] = 2'b00;
assign phi4 [24][20] = 2'b00;
assign phi4 [24][21] = 2'b10;
assign phi4 [24][22] = 2'b11;
assign phi4 [24][23] = 2'b11;
assign phi4 [25][0] = 2'b11;
assign phi4 [25][1] = 2'b00;
assign phi4 [25][2] = 2'b10;
assign phi4 [25][3] = 2'b11;
assign phi4 [25][4] = 2'b11;
assign phi4 [25][5] = 2'b10;
assign phi4 [25][6] = 2'b00;
assign phi4 [25][7] = 2'b11;
assign phi4 [25][8] = 2'b10;
assign phi4 [25][9] = 2'b11;
assign phi4 [25][10] = 2'b00;
assign phi4 [25][11] = 2'b00;
assign phi4 [25][12] = 2'b10;
assign phi4 [25][13] = 2'b00;
assign phi4 [25][14] = 2'b00;
assign phi4 [25][15] = 2'b01;
assign phi4 [25][16] = 2'b01;
assign phi4 [25][17] = 2'b01;
assign phi4 [25][18] = 2'b10;
assign phi4 [25][19] = 2'b00;
assign phi4 [25][20] = 2'b10;
assign phi4 [25][21] = 2'b00;
assign phi4 [25][22] = 2'b10;
assign phi4 [25][23] = 2'b11;
assign phi4 [26][0] = 2'b10;
assign phi4 [26][1] = 2'b01;
assign phi4 [26][2] = 2'b10;
assign phi4 [26][3] = 2'b10;
assign phi4 [26][4] = 2'b01;
assign phi4 [26][5] = 2'b01;
assign phi4 [26][6] = 2'b10;
assign phi4 [26][7] = 2'b10;
assign phi4 [26][8] = 2'b10;
assign phi4 [26][9] = 2'b01;
assign phi4 [26][10] = 2'b10;
assign phi4 [26][11] = 2'b11;
assign phi4 [26][12] = 2'b00;
assign phi4 [26][13] = 2'b01;
assign phi4 [26][14] = 2'b00;
assign phi4 [26][15] = 2'b00;
assign phi4 [26][16] = 2'b11;
assign phi4 [26][17] = 2'b11;
assign phi4 [26][18] = 2'b11;
assign phi4 [26][19] = 2'b10;
assign phi4 [26][20] = 2'b11;
assign phi4 [26][21] = 2'b10;
assign phi4 [26][22] = 2'b11;
assign phi4 [26][23] = 2'b11;
assign phi4 [27][0] = 2'b01;
assign phi4 [27][1] = 2'b11;
assign phi4 [27][2] = 2'b11;
assign phi4 [27][3] = 2'b10;
assign phi4 [27][4] = 2'b01;
assign phi4 [27][5] = 2'b01;
assign phi4 [27][6] = 2'b11;
assign phi4 [27][7] = 2'b10;
assign phi4 [27][8] = 2'b01;
assign phi4 [27][9] = 2'b00;
assign phi4 [27][10] = 2'b00;
assign phi4 [27][11] = 2'b00;
assign phi4 [27][12] = 2'b01;
assign phi4 [27][13] = 2'b10;
assign phi4 [27][14] = 2'b01;
assign phi4 [27][15] = 2'b11;
assign phi4 [27][16] = 2'b10;
assign phi4 [27][17] = 2'b01;
assign phi4 [27][18] = 2'b10;
assign phi4 [27][19] = 2'b01;
assign phi4 [27][20] = 2'b00;
assign phi4 [27][21] = 2'b10;
assign phi4 [27][22] = 2'b11;
assign phi4 [27][23] = 2'b11;
assign phi4 [28][0] = 2'b11;
assign phi4 [28][1] = 2'b00;
assign phi4 [28][2] = 2'b11;
assign phi4 [28][3] = 2'b00;
assign phi4 [28][4] = 2'b11;
assign phi4 [28][5] = 2'b00;
assign phi4 [28][6] = 2'b00;
assign phi4 [28][7] = 2'b01;
assign phi4 [28][8] = 2'b00;
assign phi4 [28][9] = 2'b11;
assign phi4 [28][10] = 2'b11;
assign phi4 [28][11] = 2'b10;
assign phi4 [28][12] = 2'b00;
assign phi4 [28][13] = 2'b01;
assign phi4 [28][14] = 2'b10;
assign phi4 [28][15] = 2'b11;
assign phi4 [28][16] = 2'b01;
assign phi4 [28][17] = 2'b00;
assign phi4 [28][18] = 2'b10;
assign phi4 [28][19] = 2'b11;
assign phi4 [28][20] = 2'b11;
assign phi4 [28][21] = 2'b11;
assign phi4 [28][22] = 2'b11;
assign phi4 [28][23] = 2'b11;
assign phi4 [29][0] = 2'b01;
assign phi4 [29][1] = 2'b11;
assign phi4 [29][2] = 2'b10;
assign phi4 [29][3] = 2'b00;
assign phi4 [29][4] = 2'b01;
assign phi4 [29][5] = 2'b10;
assign phi4 [29][6] = 2'b10;
assign phi4 [29][7] = 2'b11;
assign phi4 [29][8] = 2'b10;
assign phi4 [29][9] = 2'b01;
assign phi4 [29][10] = 2'b10;
assign phi4 [29][11] = 2'b11;
assign phi4 [29][12] = 2'b10;
assign phi4 [29][13] = 2'b11;
assign phi4 [29][14] = 2'b01;
assign phi4 [29][15] = 2'b10;
assign phi4 [29][16] = 2'b01;
assign phi4 [29][17] = 2'b00;
assign phi4 [29][18] = 2'b00;
assign phi4 [29][19] = 2'b11;
assign phi4 [29][20] = 2'b01;
assign phi4 [29][21] = 2'b11;
assign phi4 [29][22] = 2'b11;
assign phi4 [29][23] = 2'b11;

endmodule
