module phi3 (
        input   [4:0]   u,   //  Sequence number
        input   [9:0]   counter,   //  Counter of the generator
        output wire [1:0]  phi_value  //  phase of the sequence
    );

    wire [1:0] phi3 [0:29][0:17];

    assign phi_value = phi3[u][counter];
        
assign phi3 [0][0] = 2'b10;
assign phi3 [0][1] = 2'b01;
assign phi3 [0][2] = 2'b10;
assign phi3 [0][3] = 2'b11;
assign phi3 [0][4] = 2'b01;
assign phi3 [0][5] = 2'b00;
assign phi3 [0][6] = 2'b11;
assign phi3 [0][7] = 2'b10;
assign phi3 [0][8] = 2'b01;
assign phi3 [0][9] = 2'b11;
assign phi3 [0][10] = 2'b10;
assign phi3 [0][11] = 2'b10;
assign phi3 [0][12] = 2'b00;
assign phi3 [0][13] = 2'b00;
assign phi3 [0][14] = 2'b00;
assign phi3 [0][15] = 2'b10;
assign phi3 [0][16] = 2'b10;
assign phi3 [0][17] = 2'b10;
assign phi3 [1][0] = 2'b01;
assign phi3 [1][1] = 2'b11;
assign phi3 [1][2] = 2'b01;
assign phi3 [1][3] = 2'b10;
assign phi3 [1][4] = 2'b00;
assign phi3 [1][5] = 2'b01;
assign phi3 [1][6] = 2'b11;
assign phi3 [1][7] = 2'b10;
assign phi3 [1][8] = 2'b11;
assign phi3 [1][9] = 2'b11;
assign phi3 [1][10] = 2'b10;
assign phi3 [1][11] = 2'b11;
assign phi3 [1][12] = 2'b01;
assign phi3 [1][13] = 2'b00;
assign phi3 [1][14] = 2'b10;
assign phi3 [1][15] = 2'b01;
assign phi3 [1][16] = 2'b11;
assign phi3 [1][17] = 2'b01;
assign phi3 [2][0] = 2'b11;
assign phi3 [2][1] = 2'b01;
assign phi3 [2][2] = 2'b00;
assign phi3 [2][3] = 2'b10;
assign phi3 [2][4] = 2'b10;
assign phi3 [2][5] = 2'b01;
assign phi3 [2][6] = 2'b11;
assign phi3 [2][7] = 2'b10;
assign phi3 [2][8] = 2'b00;
assign phi3 [2][9] = 2'b00;
assign phi3 [2][10] = 2'b00;
assign phi3 [2][11] = 2'b00;
assign phi3 [2][12] = 2'b00;
assign phi3 [2][13] = 2'b10;
assign phi3 [2][14] = 2'b01;
assign phi3 [2][15] = 2'b10;
assign phi3 [2][16] = 2'b11;
assign phi3 [2][17] = 2'b10;
assign phi3 [3][0] = 2'b11;
assign phi3 [3][1] = 2'b11;
assign phi3 [3][2] = 2'b01;
assign phi3 [3][3] = 2'b01;
assign phi3 [3][4] = 2'b01;
assign phi3 [3][5] = 2'b00;
assign phi3 [3][6] = 2'b11;
assign phi3 [3][7] = 2'b00;
assign phi3 [3][8] = 2'b01;
assign phi3 [3][9] = 2'b01;
assign phi3 [3][10] = 2'b00;
assign phi3 [3][11] = 2'b11;
assign phi3 [3][12] = 2'b11;
assign phi3 [3][13] = 2'b01;
assign phi3 [3][14] = 2'b10;
assign phi3 [3][15] = 2'b11;
assign phi3 [3][16] = 2'b10;
assign phi3 [3][17] = 2'b00;
assign phi3 [4][0] = 2'b00;
assign phi3 [4][1] = 2'b00;
assign phi3 [4][2] = 2'b10;
assign phi3 [4][3] = 2'b10;
assign phi3 [4][4] = 2'b11;
assign phi3 [4][5] = 2'b10;
assign phi3 [4][6] = 2'b00;
assign phi3 [4][7] = 2'b11;
assign phi3 [4][8] = 2'b11;
assign phi3 [4][9] = 2'b11;
assign phi3 [4][10] = 2'b00;
assign phi3 [4][11] = 2'b11;
assign phi3 [4][12] = 2'b10;
assign phi3 [4][13] = 2'b10;
assign phi3 [4][14] = 2'b00;
assign phi3 [4][15] = 2'b10;
assign phi3 [4][16] = 2'b01;
assign phi3 [4][17] = 2'b00;
assign phi3 [5][0] = 2'b01;
assign phi3 [5][1] = 2'b11;
assign phi3 [5][2] = 2'b00;
assign phi3 [5][3] = 2'b00;
assign phi3 [5][4] = 2'b01;
assign phi3 [5][5] = 2'b10;
assign phi3 [5][6] = 2'b00;
assign phi3 [5][7] = 2'b10;
assign phi3 [5][8] = 2'b10;
assign phi3 [5][9] = 2'b11;
assign phi3 [5][10] = 2'b00;
assign phi3 [5][11] = 2'b00;
assign phi3 [5][12] = 2'b10;
assign phi3 [5][13] = 2'b01;
assign phi3 [5][14] = 2'b01;
assign phi3 [5][15] = 2'b11;
assign phi3 [5][16] = 2'b01;
assign phi3 [5][17] = 2'b10;
assign phi3 [6][0] = 2'b11;
assign phi3 [6][1] = 2'b01;
assign phi3 [6][2] = 2'b10;
assign phi3 [6][3] = 2'b00;
assign phi3 [6][4] = 2'b01;
assign phi3 [6][5] = 2'b00;
assign phi3 [6][6] = 2'b11;
assign phi3 [6][7] = 2'b10;
assign phi3 [6][8] = 2'b00;
assign phi3 [6][9] = 2'b00;
assign phi3 [6][10] = 2'b11;
assign phi3 [6][11] = 2'b00;
assign phi3 [6][12] = 2'b01;
assign phi3 [6][13] = 2'b01;
assign phi3 [6][14] = 2'b10;
assign phi3 [6][15] = 2'b11;
assign phi3 [6][16] = 2'b11;
assign phi3 [6][17] = 2'b11;
assign phi3 [7][0] = 2'b00;
assign phi3 [7][1] = 2'b00;
assign phi3 [7][2] = 2'b11;
assign phi3 [7][3] = 2'b01;
assign phi3 [7][4] = 2'b01;
assign phi3 [7][5] = 2'b00;
assign phi3 [7][6] = 2'b01;
assign phi3 [7][7] = 2'b11;
assign phi3 [7][8] = 2'b01;
assign phi3 [7][9] = 2'b10;
assign phi3 [7][10] = 2'b00;
assign phi3 [7][11] = 2'b00;
assign phi3 [7][12] = 2'b10;
assign phi3 [7][13] = 2'b00;
assign phi3 [7][14] = 2'b11;
assign phi3 [7][15] = 2'b11;
assign phi3 [7][16] = 2'b10;
assign phi3 [7][17] = 2'b01;
assign phi3 [8][0] = 2'b11;
assign phi3 [8][1] = 2'b00;
assign phi3 [8][2] = 2'b11;
assign phi3 [8][3] = 2'b11;
assign phi3 [8][4] = 2'b00;
assign phi3 [8][5] = 2'b11;
assign phi3 [8][6] = 2'b11;
assign phi3 [8][7] = 2'b01;
assign phi3 [8][8] = 2'b00;
assign phi3 [8][9] = 2'b11;
assign phi3 [8][10] = 2'b10;
assign phi3 [8][11] = 2'b11;
assign phi3 [8][12] = 2'b11;
assign phi3 [8][13] = 2'b11;
assign phi3 [8][14] = 2'b10;
assign phi3 [8][15] = 2'b00;
assign phi3 [8][16] = 2'b00;
assign phi3 [8][17] = 2'b01;
assign phi3 [9][0] = 2'b01;
assign phi3 [9][1] = 2'b10;
assign phi3 [9][2] = 2'b01;
assign phi3 [9][3] = 2'b00;
assign phi3 [9][4] = 2'b11;
assign phi3 [9][5] = 2'b11;
assign phi3 [9][6] = 2'b10;
assign phi3 [9][7] = 2'b00;
assign phi3 [9][8] = 2'b11;
assign phi3 [9][9] = 2'b11;
assign phi3 [9][10] = 2'b01;
assign phi3 [9][11] = 2'b01;
assign phi3 [9][12] = 2'b01;
assign phi3 [9][13] = 2'b00;
assign phi3 [9][14] = 2'b01;
assign phi3 [9][15] = 2'b11;
assign phi3 [9][16] = 2'b01;
assign phi3 [9][17] = 2'b11;
assign phi3 [10][0] = 2'b11;
assign phi3 [10][1] = 2'b11;
assign phi3 [10][2] = 2'b11;
assign phi3 [10][3] = 2'b00;
assign phi3 [10][4] = 2'b11;
assign phi3 [10][5] = 2'b01;
assign phi3 [10][6] = 2'b00;
assign phi3 [10][7] = 2'b00;
assign phi3 [10][8] = 2'b01;
assign phi3 [10][9] = 2'b11;
assign phi3 [10][10] = 2'b11;
assign phi3 [10][11] = 2'b00;
assign phi3 [10][12] = 2'b01;
assign phi3 [10][13] = 2'b10;
assign phi3 [10][14] = 2'b01;
assign phi3 [10][15] = 2'b11;
assign phi3 [10][16] = 2'b11;
assign phi3 [10][17] = 2'b01;
assign phi3 [11][0] = 2'b11;
assign phi3 [11][1] = 2'b11;
assign phi3 [11][2] = 2'b01;
assign phi3 [11][3] = 2'b01;
assign phi3 [11][4] = 2'b01;
assign phi3 [11][5] = 2'b10;
assign phi3 [11][6] = 2'b10;
assign phi3 [11][7] = 2'b11;
assign phi3 [11][8] = 2'b10;
assign phi3 [11][9] = 2'b10;
assign phi3 [11][10] = 2'b10;
assign phi3 [11][11] = 2'b01;
assign phi3 [11][12] = 2'b00;
assign phi3 [11][13] = 2'b11;
assign phi3 [11][14] = 2'b11;
assign phi3 [11][15] = 2'b10;
assign phi3 [11][16] = 2'b01;
assign phi3 [11][17] = 2'b10;
assign phi3 [12][0] = 2'b11;
assign phi3 [12][1] = 2'b10;
assign phi3 [12][2] = 2'b11;
assign phi3 [12][3] = 2'b11;
assign phi3 [12][4] = 2'b00;
assign phi3 [12][5] = 2'b00;
assign phi3 [12][6] = 2'b10;
assign phi3 [12][7] = 2'b11;
assign phi3 [12][8] = 2'b10;
assign phi3 [12][9] = 2'b11;
assign phi3 [12][10] = 2'b10;
assign phi3 [12][11] = 2'b10;
assign phi3 [12][12] = 2'b01;
assign phi3 [12][13] = 2'b01;
assign phi3 [12][14] = 2'b10;
assign phi3 [12][15] = 2'b01;
assign phi3 [12][16] = 2'b00;
assign phi3 [12][17] = 2'b01;
assign phi3 [13][0] = 2'b00;
assign phi3 [13][1] = 2'b00;
assign phi3 [13][2] = 2'b11;
assign phi3 [13][3] = 2'b11;
assign phi3 [13][4] = 2'b11;
assign phi3 [13][5] = 2'b11;
assign phi3 [13][6] = 2'b00;
assign phi3 [13][7] = 2'b01;
assign phi3 [13][8] = 2'b11;
assign phi3 [13][9] = 2'b01;
assign phi3 [13][10] = 2'b01;
assign phi3 [13][11] = 2'b00;
assign phi3 [13][12] = 2'b11;
assign phi3 [13][13] = 2'b10;
assign phi3 [13][14] = 2'b01;
assign phi3 [13][15] = 2'b10;
assign phi3 [13][16] = 2'b11;
assign phi3 [13][17] = 2'b00;
assign phi3 [14][0] = 2'b11;
assign phi3 [14][1] = 2'b01;
assign phi3 [14][2] = 2'b10;
assign phi3 [14][3] = 2'b11;
assign phi3 [14][4] = 2'b10;
assign phi3 [14][5] = 2'b11;
assign phi3 [14][6] = 2'b00;
assign phi3 [14][7] = 2'b00;
assign phi3 [14][8] = 2'b11;
assign phi3 [14][9] = 2'b11;
assign phi3 [14][10] = 2'b10;
assign phi3 [14][11] = 2'b10;
assign phi3 [14][12] = 2'b01;
assign phi3 [14][13] = 2'b11;
assign phi3 [14][14] = 2'b00;
assign phi3 [14][15] = 2'b01;
assign phi3 [14][16] = 2'b00;
assign phi3 [14][17] = 2'b00;
assign phi3 [15][0] = 2'b01;
assign phi3 [15][1] = 2'b00;
assign phi3 [15][2] = 2'b11;
assign phi3 [15][3] = 2'b00;
assign phi3 [15][4] = 2'b11;
assign phi3 [15][5] = 2'b01;
assign phi3 [15][6] = 2'b01;
assign phi3 [15][7] = 2'b10;
assign phi3 [15][8] = 2'b11;
assign phi3 [15][9] = 2'b11;
assign phi3 [15][10] = 2'b10;
assign phi3 [15][11] = 2'b11;
assign phi3 [15][12] = 2'b11;
assign phi3 [15][13] = 2'b01;
assign phi3 [15][14] = 2'b11;
assign phi3 [15][15] = 2'b10;
assign phi3 [15][16] = 2'b00;
assign phi3 [15][17] = 2'b01;
assign phi3 [16][0] = 2'b11;
assign phi3 [16][1] = 2'b10;
assign phi3 [16][2] = 2'b11;
assign phi3 [16][3] = 2'b10;
assign phi3 [16][4] = 2'b11;
assign phi3 [16][5] = 2'b00;
assign phi3 [16][6] = 2'b01;
assign phi3 [16][7] = 2'b11;
assign phi3 [16][8] = 2'b10;
assign phi3 [16][9] = 2'b01;
assign phi3 [16][10] = 2'b01;
assign phi3 [16][11] = 2'b01;
assign phi3 [16][12] = 2'b00;
assign phi3 [16][13] = 2'b10;
assign phi3 [16][14] = 2'b11;
assign phi3 [16][15] = 2'b01;
assign phi3 [16][16] = 2'b10;
assign phi3 [16][17] = 2'b11;
assign phi3 [17][0] = 2'b11;
assign phi3 [17][1] = 2'b10;
assign phi3 [17][2] = 2'b01;
assign phi3 [17][3] = 2'b01;
assign phi3 [17][4] = 2'b10;
assign phi3 [17][5] = 2'b01;
assign phi3 [17][6] = 2'b10;
assign phi3 [17][7] = 2'b11;
assign phi3 [17][8] = 2'b10;
assign phi3 [17][9] = 2'b00;
assign phi3 [17][10] = 2'b10;
assign phi3 [17][11] = 2'b11;
assign phi3 [17][12] = 2'b10;
assign phi3 [17][13] = 2'b10;
assign phi3 [17][14] = 2'b10;
assign phi3 [17][15] = 2'b01;
assign phi3 [17][16] = 2'b01;
assign phi3 [17][17] = 2'b00;
assign phi3 [18][0] = 2'b11;
assign phi3 [18][1] = 2'b00;
assign phi3 [18][2] = 2'b11;
assign phi3 [18][3] = 2'b10;
assign phi3 [18][4] = 2'b10;
assign phi3 [18][5] = 2'b01;
assign phi3 [18][6] = 2'b00;
assign phi3 [18][7] = 2'b11;
assign phi3 [18][8] = 2'b11;
assign phi3 [18][9] = 2'b11;
assign phi3 [18][10] = 2'b10;
assign phi3 [18][11] = 2'b11;
assign phi3 [18][12] = 2'b11;
assign phi3 [18][13] = 2'b00;
assign phi3 [18][14] = 2'b00;
assign phi3 [18][15] = 2'b00;
assign phi3 [18][16] = 2'b10;
assign phi3 [18][17] = 2'b10;
assign phi3 [19][0] = 2'b01;
assign phi3 [19][1] = 2'b01;
assign phi3 [19][2] = 2'b01;
assign phi3 [19][3] = 2'b11;
assign phi3 [19][4] = 2'b10;
assign phi3 [19][5] = 2'b11;
assign phi3 [19][6] = 2'b10;
assign phi3 [19][7] = 2'b01;
assign phi3 [19][8] = 2'b10;
assign phi3 [19][9] = 2'b00;
assign phi3 [19][10] = 2'b10;
assign phi3 [19][11] = 2'b11;
assign phi3 [19][12] = 2'b00;
assign phi3 [19][13] = 2'b11;
assign phi3 [19][14] = 2'b11;
assign phi3 [19][15] = 2'b10;
assign phi3 [19][16] = 2'b01;
assign phi3 [19][17] = 2'b01;
assign phi3 [20][0] = 2'b11;
assign phi3 [20][1] = 2'b00;
assign phi3 [20][2] = 2'b00;
assign phi3 [20][3] = 2'b11;
assign phi3 [20][4] = 2'b00;
assign phi3 [20][5] = 2'b00;
assign phi3 [20][6] = 2'b01;
assign phi3 [20][7] = 2'b11;
assign phi3 [20][8] = 2'b10;
assign phi3 [20][9] = 2'b11;
assign phi3 [20][10] = 2'b10;
assign phi3 [20][11] = 2'b01;
assign phi3 [20][12] = 2'b11;
assign phi3 [20][13] = 2'b01;
assign phi3 [20][14] = 2'b10;
assign phi3 [20][15] = 2'b10;
assign phi3 [20][16] = 2'b10;
assign phi3 [20][17] = 2'b11;
assign phi3 [21][0] = 2'b00;
assign phi3 [21][1] = 2'b11;
assign phi3 [21][2] = 2'b10;
assign phi3 [21][3] = 2'b11;
assign phi3 [21][4] = 2'b01;
assign phi3 [21][5] = 2'b01;
assign phi3 [21][6] = 2'b10;
assign phi3 [21][7] = 2'b11;
assign phi3 [21][8] = 2'b00;
assign phi3 [21][9] = 2'b11;
assign phi3 [21][10] = 2'b11;
assign phi3 [21][11] = 2'b10;
assign phi3 [21][12] = 2'b11;
assign phi3 [21][13] = 2'b10;
assign phi3 [21][14] = 2'b00;
assign phi3 [21][15] = 2'b01;
assign phi3 [21][16] = 2'b01;
assign phi3 [21][17] = 2'b01;
assign phi3 [22][0] = 2'b11;
assign phi3 [22][1] = 2'b11;
assign phi3 [22][2] = 2'b00;
assign phi3 [22][3] = 2'b10;
assign phi3 [22][4] = 2'b10;
assign phi3 [22][5] = 2'b00;
assign phi3 [22][6] = 2'b00;
assign phi3 [22][7] = 2'b11;
assign phi3 [22][8] = 2'b10;
assign phi3 [22][9] = 2'b01;
assign phi3 [22][10] = 2'b01;
assign phi3 [22][11] = 2'b01;
assign phi3 [22][12] = 2'b01;
assign phi3 [22][13] = 2'b10;
assign phi3 [22][14] = 2'b01;
assign phi3 [22][15] = 2'b00;
assign phi3 [22][16] = 2'b01;
assign phi3 [22][17] = 2'b00;
assign phi3 [23][0] = 2'b01;
assign phi3 [23][1] = 2'b10;
assign phi3 [23][2] = 2'b11;
assign phi3 [23][3] = 2'b00;
assign phi3 [23][4] = 2'b11;
assign phi3 [23][5] = 2'b11;
assign phi3 [23][6] = 2'b11;
assign phi3 [23][7] = 2'b01;
assign phi3 [23][8] = 2'b01;
assign phi3 [23][9] = 2'b10;
assign phi3 [23][10] = 2'b00;
assign phi3 [23][11] = 2'b11;
assign phi3 [23][12] = 2'b10;
assign phi3 [23][13] = 2'b01;
assign phi3 [23][14] = 2'b00;
assign phi3 [23][15] = 2'b00;
assign phi3 [23][16] = 2'b01;
assign phi3 [23][17] = 2'b01;
assign phi3 [24][0] = 2'b01;
assign phi3 [24][1] = 2'b10;
assign phi3 [24][2] = 2'b10;
assign phi3 [24][3] = 2'b00;
assign phi3 [24][4] = 2'b11;
assign phi3 [24][5] = 2'b10;
assign phi3 [24][6] = 2'b11;
assign phi3 [24][7] = 2'b10;
assign phi3 [24][8] = 2'b11;
assign phi3 [24][9] = 2'b11;
assign phi3 [24][10] = 2'b10;
assign phi3 [24][11] = 2'b11;
assign phi3 [24][12] = 2'b00;
assign phi3 [24][13] = 2'b00;
assign phi3 [24][14] = 2'b00;
assign phi3 [24][15] = 2'b11;
assign phi3 [24][16] = 2'b11;
assign phi3 [24][17] = 2'b01;
assign phi3 [25][0] = 2'b11;
assign phi3 [25][1] = 2'b11;
assign phi3 [25][2] = 2'b00;
assign phi3 [25][3] = 2'b11;
assign phi3 [25][4] = 2'b01;
assign phi3 [25][5] = 2'b01;
assign phi3 [25][6] = 2'b01;
assign phi3 [25][7] = 2'b10;
assign phi3 [25][8] = 2'b01;
assign phi3 [25][9] = 2'b00;
assign phi3 [25][10] = 2'b00;
assign phi3 [25][11] = 2'b11;
assign phi3 [25][12] = 2'b11;
assign phi3 [25][13] = 2'b11;
assign phi3 [25][14] = 2'b01;
assign phi3 [25][15] = 2'b11;
assign phi3 [25][16] = 2'b10;
assign phi3 [25][17] = 2'b10;
assign phi3 [26][0] = 2'b11;
assign phi3 [26][1] = 2'b10;
assign phi3 [26][2] = 2'b10;
assign phi3 [26][3] = 2'b11;
assign phi3 [26][4] = 2'b00;
assign phi3 [26][5] = 2'b11;
assign phi3 [26][6] = 2'b01;
assign phi3 [26][7] = 2'b10;
assign phi3 [26][8] = 2'b10;
assign phi3 [26][9] = 2'b11;
assign phi3 [26][10] = 2'b01;
assign phi3 [26][11] = 2'b01;
assign phi3 [26][12] = 2'b11;
assign phi3 [26][13] = 2'b10;
assign phi3 [26][14] = 2'b01;
assign phi3 [26][15] = 2'b10;
assign phi3 [26][16] = 2'b10;
assign phi3 [26][17] = 2'b10;
assign phi3 [27][0] = 2'b11;
assign phi3 [27][1] = 2'b11;
assign phi3 [27][2] = 2'b01;
assign phi3 [27][3] = 2'b01;
assign phi3 [27][4] = 2'b11;
assign phi3 [27][5] = 2'b00;
assign phi3 [27][6] = 2'b01;
assign phi3 [27][7] = 2'b10;
assign phi3 [27][8] = 2'b11;
assign phi3 [27][9] = 2'b00;
assign phi3 [27][10] = 2'b10;
assign phi3 [27][11] = 2'b11;
assign phi3 [27][12] = 2'b01;
assign phi3 [27][13] = 2'b11;
assign phi3 [27][14] = 2'b10;
assign phi3 [27][15] = 2'b10;
assign phi3 [27][16] = 2'b10;
assign phi3 [27][17] = 2'b01;
assign phi3 [28][0] = 2'b10;
assign phi3 [28][1] = 2'b11;
assign phi3 [28][2] = 2'b00;
assign phi3 [28][3] = 2'b11;
assign phi3 [28][4] = 2'b11;
assign phi3 [28][5] = 2'b11;
assign phi3 [28][6] = 2'b00;
assign phi3 [28][7] = 2'b00;
assign phi3 [28][8] = 2'b01;
assign phi3 [28][9] = 2'b01;
assign phi3 [28][10] = 2'b11;
assign phi3 [28][11] = 2'b01;
assign phi3 [28][12] = 2'b01;
assign phi3 [28][13] = 2'b11;
assign phi3 [28][14] = 2'b10;
assign phi3 [28][15] = 2'b01;
assign phi3 [28][16] = 2'b11;
assign phi3 [28][17] = 2'b00;
assign phi3 [29][0] = 2'b11;
assign phi3 [29][1] = 2'b01;
assign phi3 [29][2] = 2'b00;
assign phi3 [29][3] = 2'b10;
assign phi3 [29][4] = 2'b10;
assign phi3 [29][5] = 2'b10;
assign phi3 [29][6] = 2'b10;
assign phi3 [29][7] = 2'b00;
assign phi3 [29][8] = 2'b10;
assign phi3 [29][9] = 2'b01;
assign phi3 [29][10] = 2'b01;
assign phi3 [29][11] = 2'b11;
assign phi3 [29][12] = 2'b10;
assign phi3 [29][13] = 2'b00;
assign phi3 [29][14] = 2'b01;
assign phi3 [29][15] = 2'b10;
assign phi3 [29][16] = 2'b01;
assign phi3 [29][17] = 2'b10;

endmodule
