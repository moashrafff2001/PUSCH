module phi1 (
        input   [4:0]   u,   //  Sequence number
        input   [9:0]   counter,   //  Counter of the generator
        output  [1:0]  phi_value  //  phase of the sequence
    );

    wire [1:0] phi1 [0:29][0:5];
    assign phi_value = phi1[u][counter];
assign phi1 [0][0] = 2'b11;
assign phi1 [0][1] = 2'b10;
assign phi1 [0][2] = 2'b01;
assign phi1 [0][3] = 2'b01;
assign phi1 [0][4] = 2'b10;
assign phi1 [0][5] = 2'b11;
assign phi1 [1][0] = 2'b11;
assign phi1 [1][1] = 2'b01;
assign phi1 [1][2] = 2'b10;
assign phi1 [1][3] = 2'b10;
assign phi1 [1][4] = 2'b01;
assign phi1 [1][5] = 2'b11;
assign phi1 [2][0] = 2'b11;
assign phi1 [2][1] = 2'b11;
assign phi1 [2][2] = 2'b11;
assign phi1 [2][3] = 2'b01;
assign phi1 [2][4] = 2'b00;
assign phi1 [2][5] = 2'b11;
assign phi1 [3][0] = 2'b00;
assign phi1 [3][1] = 2'b00;
assign phi1 [3][2] = 2'b00;
assign phi1 [3][3] = 2'b01;
assign phi1 [3][4] = 2'b10;
assign phi1 [3][5] = 2'b11;
assign phi1 [4][0] = 2'b00;
assign phi1 [4][1] = 2'b00;
assign phi1 [4][2] = 2'b00;
assign phi1 [4][3] = 2'b11;
assign phi1 [4][4] = 2'b10;
assign phi1 [4][5] = 2'b01;
assign phi1 [5][0] = 2'b11;
assign phi1 [5][1] = 2'b00;
assign phi1 [5][2] = 2'b10;
assign phi1 [5][3] = 2'b11;
assign phi1 [5][4] = 2'b11;
assign phi1 [5][5] = 2'b11;
assign phi1 [6][0] = 2'b11;
assign phi1 [6][1] = 2'b00;
assign phi1 [6][2] = 2'b01;
assign phi1 [6][3] = 2'b11;
assign phi1 [6][4] = 2'b11;
assign phi1 [6][5] = 2'b11;
assign phi1 [7][0] = 2'b11;
assign phi1 [7][1] = 2'b10;
assign phi1 [7][2] = 2'b00;
assign phi1 [7][3] = 2'b11;
assign phi1 [7][4] = 2'b00;
assign phi1 [7][5] = 2'b10;
assign phi1 [8][0] = 2'b11;
assign phi1 [8][1] = 2'b10;
assign phi1 [8][2] = 2'b11;
assign phi1 [8][3] = 2'b00;
assign phi1 [8][4] = 2'b11;
assign phi1 [8][5] = 2'b11;
assign phi1 [9][0] = 2'b11;
assign phi1 [9][1] = 2'b11;
assign phi1 [9][2] = 2'b00;
assign phi1 [9][3] = 2'b11;
assign phi1 [9][4] = 2'b01;
assign phi1 [9][5] = 2'b11;
assign phi1 [10][0] = 2'b11;
assign phi1 [10][1] = 2'b00;
assign phi1 [10][2] = 2'b01;
assign phi1 [10][3] = 2'b00;
assign phi1 [10][4] = 2'b11;
assign phi1 [10][5] = 2'b11;
assign phi1 [11][0] = 2'b11;
assign phi1 [11][1] = 2'b10;
assign phi1 [11][2] = 2'b11;
assign phi1 [11][3] = 2'b00;
assign phi1 [11][4] = 2'b00;
assign phi1 [11][5] = 2'b11;
assign phi1 [12][0] = 2'b00;
assign phi1 [12][1] = 2'b00;
assign phi1 [12][2] = 2'b01;
assign phi1 [12][3] = 2'b10;
assign phi1 [12][4] = 2'b11;
assign phi1 [12][5] = 2'b01;
assign phi1 [13][0] = 2'b00;
assign phi1 [13][1] = 2'b00;
assign phi1 [13][2] = 2'b01;
assign phi1 [13][3] = 2'b01;
assign phi1 [13][4] = 2'b10;
assign phi1 [13][5] = 2'b01;
assign phi1 [14][0] = 2'b00;
assign phi1 [14][1] = 2'b00;
assign phi1 [14][2] = 2'b00;
assign phi1 [14][3] = 2'b11;
assign phi1 [14][4] = 2'b01;
assign phi1 [14][5] = 2'b10;
assign phi1 [15][0] = 2'b00;
assign phi1 [15][1] = 2'b00;
assign phi1 [15][2] = 2'b00;
assign phi1 [15][3] = 2'b10;
assign phi1 [15][4] = 2'b01;
assign phi1 [15][5] = 2'b11;
assign phi1 [16][0] = 2'b11;
assign phi1 [16][1] = 2'b10;
assign phi1 [16][2] = 2'b10;
assign phi1 [16][3] = 2'b10;
assign phi1 [16][4] = 2'b01;
assign phi1 [16][5] = 2'b10;
assign phi1 [17][0] = 2'b11;
assign phi1 [17][1] = 2'b11;
assign phi1 [17][2] = 2'b10;
assign phi1 [17][3] = 2'b00;
assign phi1 [17][4] = 2'b10;
assign phi1 [17][5] = 2'b11;
assign phi1 [18][0] = 2'b11;
assign phi1 [18][1] = 2'b11;
assign phi1 [18][2] = 2'b11;
assign phi1 [18][3] = 2'b00;
assign phi1 [18][4] = 2'b11;
assign phi1 [18][5] = 2'b10;
assign phi1 [19][0] = 2'b11;
assign phi1 [19][1] = 2'b00;
assign phi1 [19][2] = 2'b00;
assign phi1 [19][3] = 2'b11;
assign phi1 [19][4] = 2'b10;
assign phi1 [19][5] = 2'b11;
assign phi1 [20][0] = 2'b11;
assign phi1 [20][1] = 2'b01;
assign phi1 [20][2] = 2'b11;
assign phi1 [20][3] = 2'b00;
assign phi1 [20][4] = 2'b00;
assign phi1 [20][5] = 2'b11;
assign phi1 [21][0] = 2'b11;
assign phi1 [21][1] = 2'b00;
assign phi1 [21][2] = 2'b11;
assign phi1 [21][3] = 2'b11;
assign phi1 [21][4] = 2'b11;
assign phi1 [21][5] = 2'b10;
assign phi1 [22][0] = 2'b00;
assign phi1 [22][1] = 2'b00;
assign phi1 [22][2] = 2'b11;
assign phi1 [22][3] = 2'b01;
assign phi1 [22][4] = 2'b00;
assign phi1 [22][5] = 2'b01;
assign phi1 [23][0] = 2'b00;
assign phi1 [23][1] = 2'b00;
assign phi1 [23][2] = 2'b11;
assign phi1 [23][3] = 2'b11;
assign phi1 [23][4] = 2'b00;
assign phi1 [23][5] = 2'b11;
assign phi1 [24][0] = 2'b00;
assign phi1 [24][1] = 2'b00;
assign phi1 [24][2] = 2'b01;
assign phi1 [24][3] = 2'b10;
assign phi1 [24][4] = 2'b01;
assign phi1 [24][5] = 2'b01;
assign phi1 [25][0] = 2'b00;
assign phi1 [25][1] = 2'b00;
assign phi1 [25][2] = 2'b11;
assign phi1 [25][3] = 2'b00;
assign phi1 [25][4] = 2'b01;
assign phi1 [25][5] = 2'b01;
assign phi1 [26][0] = 2'b00;
assign phi1 [26][1] = 2'b00;
assign phi1 [26][2] = 2'b10;
assign phi1 [26][3] = 2'b10;
assign phi1 [26][4] = 2'b01;
assign phi1 [26][5] = 2'b10;
assign phi1 [27][0] = 2'b00;
assign phi1 [27][1] = 2'b00;
assign phi1 [27][2] = 2'b10;
assign phi1 [27][3] = 2'b01;
assign phi1 [27][4] = 2'b10;
assign phi1 [27][5] = 2'b10;
assign phi1 [28][0] = 2'b00;
assign phi1 [28][1] = 2'b00;
assign phi1 [28][2] = 2'b10;
assign phi1 [28][3] = 2'b01;
assign phi1 [28][4] = 2'b11;
assign phi1 [28][5] = 2'b10;
assign phi1 [29][0] = 2'b00;
assign phi1 [29][1] = 2'b00;
assign phi1 [29][2] = 2'b11;
assign phi1 [29][3] = 2'b00;
assign phi1 [29][4] = 2'b10;
assign phi1 [29][5] = 2'b10;

endmodule
